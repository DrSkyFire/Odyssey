//=============================================================================
// 文件名: char_rom_16x32.v
// 描述: 16x32点阵字符ROM - 支持0-9数字及常用字符
// 美观的大字体设计，适合HDMI显示
//=============================================================================

module char_rom_16x32 (
    input  wire [5:0]   char_code,      // 字符编码
    input  wire [4:0]   row,            // 行号 (0-31)
    output reg  [15:0]  pixel_row       // 16位像素行数据
);

always @(*) begin
    case (char_code)
        //=====================================================
        // '0' - ASCII 48
        //=====================================================
        6'd0: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0001111111111000;
                5'd2:  pixel_row = 16'b0011111111111100;
                5'd3:  pixel_row = 16'b0111110000111110;
                5'd4:  pixel_row = 16'b0111100000011110;
                5'd5:  pixel_row = 16'b1111000000001111;
                5'd6:  pixel_row = 16'b1111000000001111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1110000000000111;
                5'd9:  pixel_row = 16'b1110000000000111;
                5'd10: pixel_row = 16'b1110000000000111;
                5'd11: pixel_row = 16'b1110000000000111;
                5'd12: pixel_row = 16'b1110000000000111;
                5'd13: pixel_row = 16'b1110000000000111;
                5'd14: pixel_row = 16'b1110000000000111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                5'd17: pixel_row = 16'b1110000000000111;
                5'd18: pixel_row = 16'b1110000000000111;
                5'd19: pixel_row = 16'b1110000000000111;
                5'd20: pixel_row = 16'b1110000000000111;
                5'd21: pixel_row = 16'b1110000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1110000000000111;
                5'd24: pixel_row = 16'b1111000000001111;
                5'd25: pixel_row = 16'b1111000000001111;
                5'd26: pixel_row = 16'b0111100000011110;
                5'd27: pixel_row = 16'b0111110000111110;
                5'd28: pixel_row = 16'b0011111111111100;
                5'd29: pixel_row = 16'b0001111111111000;
                5'd30: pixel_row = 16'b0000111111110000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '1' - ASCII 49
        //=====================================================
        6'd1: begin
            case (row)
                5'd0:  pixel_row = 16'b0000001110000000;
                5'd1:  pixel_row = 16'b0000011110000000;
                5'd2:  pixel_row = 16'b0000111110000000;
                5'd3:  pixel_row = 16'b0001111110000000;
                5'd4:  pixel_row = 16'b0011111110000000;
                5'd5:  pixel_row = 16'b0011100110000000;
                5'd6:  pixel_row = 16'b0000000110000000;
                5'd7:  pixel_row = 16'b0000000110000000;
                5'd8:  pixel_row = 16'b0000000110000000;
                5'd9:  pixel_row = 16'b0000000110000000;
                5'd10: pixel_row = 16'b0000000110000000;
                5'd11: pixel_row = 16'b0000000110000000;
                5'd12: pixel_row = 16'b0000000110000000;
                5'd13: pixel_row = 16'b0000000110000000;
                5'd14: pixel_row = 16'b0000000110000000;
                5'd15: pixel_row = 16'b0000000110000000;
                5'd16: pixel_row = 16'b0000000110000000;
                5'd17: pixel_row = 16'b0000000110000000;
                5'd18: pixel_row = 16'b0000000110000000;
                5'd19: pixel_row = 16'b0000000110000000;
                5'd20: pixel_row = 16'b0000000110000000;
                5'd21: pixel_row = 16'b0000000110000000;
                5'd22: pixel_row = 16'b0000000110000000;
                5'd23: pixel_row = 16'b0000000110000000;
                5'd24: pixel_row = 16'b0000000110000000;
                5'd25: pixel_row = 16'b0000000110000000;
                5'd26: pixel_row = 16'b0000000110000000;
                5'd27: pixel_row = 16'b0111111111111110;
                5'd28: pixel_row = 16'b0111111111111110;
                5'd29: pixel_row = 16'b0111111111111110;
                5'd30: pixel_row = 16'b0111111111111110;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '2' - ASCII 50
        //=====================================================
        6'd2: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0011111111111100;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111100000011110;
                5'd4:  pixel_row = 16'b1110000000001111;
                5'd5:  pixel_row = 16'b1110000000000111;
                5'd6:  pixel_row = 16'b0000000000000111;
                5'd7:  pixel_row = 16'b0000000000000111;
                5'd8:  pixel_row = 16'b0000000000001111;
                5'd9:  pixel_row = 16'b0000000000011110;
                5'd10: pixel_row = 16'b0000000000111100;
                5'd11: pixel_row = 16'b0000000001111000;
                5'd12: pixel_row = 16'b0000000011110000;
                5'd13: pixel_row = 16'b0000000111100000;
                5'd14: pixel_row = 16'b0000001111000000;
                5'd15: pixel_row = 16'b0000011110000000;
                5'd16: pixel_row = 16'b0000111100000000;
                5'd17: pixel_row = 16'b0001111000000000;
                5'd18: pixel_row = 16'b0011110000000000;
                5'd19: pixel_row = 16'b0111100000000000;
                5'd20: pixel_row = 16'b0111000000000000;
                5'd21: pixel_row = 16'b1110000000000000;
                5'd22: pixel_row = 16'b1110000000000000;
                5'd23: pixel_row = 16'b1110000000000000;
                5'd24: pixel_row = 16'b1110000000000000;
                5'd25: pixel_row = 16'b1111000000000000;
                5'd26: pixel_row = 16'b1111111111111111;
                5'd27: pixel_row = 16'b1111111111111111;
                5'd28: pixel_row = 16'b1111111111111111;
                5'd29: pixel_row = 16'b1111111111111111;
                5'd30: pixel_row = 16'b1111111111111111;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '3' - ASCII 51
        //=====================================================
        6'd3: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0011111111111100;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111000000011110;
                5'd4:  pixel_row = 16'b1110000000001111;
                5'd5:  pixel_row = 16'b0000000000000111;
                5'd6:  pixel_row = 16'b0000000000000111;
                5'd7:  pixel_row = 16'b0000000000001110;
                5'd8:  pixel_row = 16'b0000000000111100;
                5'd9:  pixel_row = 16'b0000000111111000;
                5'd10: pixel_row = 16'b0000000111111000;
                5'd11: pixel_row = 16'b0000000111111000;
                5'd12: pixel_row = 16'b0000000111111000;
                5'd13: pixel_row = 16'b0000000111111000;
                5'd14: pixel_row = 16'b0000000000111100;
                5'd15: pixel_row = 16'b0000000000001110;
                5'd16: pixel_row = 16'b0000000000000111;
                5'd17: pixel_row = 16'b0000000000000111;
                5'd18: pixel_row = 16'b0000000000000111;
                5'd19: pixel_row = 16'b0000000000000111;
                5'd20: pixel_row = 16'b0000000000000111;
                5'd21: pixel_row = 16'b0000000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1110000000001111;
                5'd24: pixel_row = 16'b1111000000001111;
                5'd25: pixel_row = 16'b0111100000011110;
                5'd26: pixel_row = 16'b0111110000111110;
                5'd27: pixel_row = 16'b0011111111111100;
                5'd28: pixel_row = 16'b0001111111111000;
                5'd29: pixel_row = 16'b0000111111110000;
                5'd30: pixel_row = 16'b0000011111100000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '4' - ASCII 52
        //=====================================================
        6'd4: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000001111000;
                5'd1:  pixel_row = 16'b0000000011111000;
                5'd2:  pixel_row = 16'b0000000111111000;
                5'd3:  pixel_row = 16'b0000000111011000;
                5'd4:  pixel_row = 16'b0000001110011000;
                5'd5:  pixel_row = 16'b0000011100011000;
                5'd6:  pixel_row = 16'b0000011100011000;
                5'd7:  pixel_row = 16'b0000111000011000;
                5'd8:  pixel_row = 16'b0001110000011000;
                5'd9:  pixel_row = 16'b0011100000011000;
                5'd10: pixel_row = 16'b0011100000011000;
                5'd11: pixel_row = 16'b0111000000011000;
                5'd12: pixel_row = 16'b1110000000011000;
                5'd13: pixel_row = 16'b1110000000011000;
                5'd14: pixel_row = 16'b1100000000011000;
                5'd15: pixel_row = 16'b1111111111111111;
                5'd16: pixel_row = 16'b1111111111111111;
                5'd17: pixel_row = 16'b1111111111111111;
                5'd18: pixel_row = 16'b0000000000011000;
                5'd19: pixel_row = 16'b0000000000011000;
                5'd20: pixel_row = 16'b0000000000011000;
                5'd21: pixel_row = 16'b0000000000011000;
                5'd22: pixel_row = 16'b0000000000011000;
                5'd23: pixel_row = 16'b0000000000011000;
                5'd24: pixel_row = 16'b0000000000011000;
                5'd25: pixel_row = 16'b0000000000011000;
                5'd26: pixel_row = 16'b0000000000011000;
                5'd27: pixel_row = 16'b0000000000011000;
                5'd28: pixel_row = 16'b0000000000011000;
                5'd29: pixel_row = 16'b0000000000011000;
                5'd30: pixel_row = 16'b0000000000011000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '5' - ASCII 53
        //=====================================================
        6'd5: begin
            case (row)
                5'd0:  pixel_row = 16'b0111111111111110;
                5'd1:  pixel_row = 16'b0111111111111110;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111000000000000;
                5'd4:  pixel_row = 16'b0111000000000000;
                5'd5:  pixel_row = 16'b1110000000000000;
                5'd6:  pixel_row = 16'b1110000000000000;
                5'd7:  pixel_row = 16'b1110000000000000;
                5'd8:  pixel_row = 16'b1110111111100000;
                5'd9:  pixel_row = 16'b1111111111111000;
                5'd10: pixel_row = 16'b1111111111111100;
                5'd11: pixel_row = 16'b1111100000111110;
                5'd12: pixel_row = 16'b1110000000011110;
                5'd13: pixel_row = 16'b0000000000001111;
                5'd14: pixel_row = 16'b0000000000000111;
                5'd15: pixel_row = 16'b0000000000000111;
                5'd16: pixel_row = 16'b0000000000000111;
                5'd17: pixel_row = 16'b0000000000000111;
                5'd18: pixel_row = 16'b0000000000000111;
                5'd19: pixel_row = 16'b0000000000000111;
                5'd20: pixel_row = 16'b0000000000000111;
                5'd21: pixel_row = 16'b0000000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1110000000001111;
                5'd24: pixel_row = 16'b1111000000001111;
                5'd25: pixel_row = 16'b0111100000011110;
                5'd26: pixel_row = 16'b0111110000111110;
                5'd27: pixel_row = 16'b0011111111111100;
                5'd28: pixel_row = 16'b0001111111111000;
                5'd29: pixel_row = 16'b0000111111110000;
                5'd30: pixel_row = 16'b0000011111100000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '6' - ASCII 54
        //=====================================================
        6'd6: begin
            case (row)
                5'd0:  pixel_row = 16'b0000011111110000;
                5'd1:  pixel_row = 16'b0001111111111000;
                5'd2:  pixel_row = 16'b0011111111111100;
                5'd3:  pixel_row = 16'b0111110000000000;
                5'd4:  pixel_row = 16'b0111100000000000;
                5'd5:  pixel_row = 16'b1111000000000000;
                5'd6:  pixel_row = 16'b1110000000000000;
                5'd7:  pixel_row = 16'b1110000000000000;
                5'd8:  pixel_row = 16'b1110011111100000;
                5'd9:  pixel_row = 16'b1110111111111000;
                5'd10: pixel_row = 16'b1111111111111100;
                5'd11: pixel_row = 16'b1111110000111110;
                5'd12: pixel_row = 16'b1111100000011110;
                5'd13: pixel_row = 16'b1111000000001111;
                5'd14: pixel_row = 16'b1110000000000111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                5'd17: pixel_row = 16'b1110000000000111;
                5'd18: pixel_row = 16'b1110000000000111;
                5'd19: pixel_row = 16'b1110000000000111;
                5'd20: pixel_row = 16'b1110000000000111;
                5'd21: pixel_row = 16'b1110000000000111;
                5'd22: pixel_row = 16'b1110000000001111;
                5'd23: pixel_row = 16'b1111000000001111;
                5'd24: pixel_row = 16'b0111100000011110;
                5'd25: pixel_row = 16'b0111110000111110;
                5'd26: pixel_row = 16'b0011111111111100;
                5'd27: pixel_row = 16'b0001111111111000;
                5'd28: pixel_row = 16'b0000111111110000;
                5'd29: pixel_row = 16'b0000011111100000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '7' - ASCII 55
        //=====================================================
        6'd7: begin
            case (row)
                5'd0:  pixel_row = 16'b1111111111111111;
                5'd1:  pixel_row = 16'b1111111111111111;
                5'd2:  pixel_row = 16'b1111111111111111;
                5'd3:  pixel_row = 16'b1111111111111111;
                5'd4:  pixel_row = 16'b0000000000000111;
                5'd5:  pixel_row = 16'b0000000000001110;
                5'd6:  pixel_row = 16'b0000000000011100;
                5'd7:  pixel_row = 16'b0000000000111000;
                5'd8:  pixel_row = 16'b0000000000111000;
                5'd9:  pixel_row = 16'b0000000001110000;
                5'd10: pixel_row = 16'b0000000011100000;
                5'd11: pixel_row = 16'b0000000011100000;
                5'd12: pixel_row = 16'b0000000111000000;
                5'd13: pixel_row = 16'b0000000111000000;
                5'd14: pixel_row = 16'b0000001110000000;
                5'd15: pixel_row = 16'b0000001110000000;
                5'd16: pixel_row = 16'b0000011100000000;
                5'd17: pixel_row = 16'b0000011100000000;
                5'd18: pixel_row = 16'b0000111000000000;
                5'd19: pixel_row = 16'b0000111000000000;
                5'd20: pixel_row = 16'b0001110000000000;
                5'd21: pixel_row = 16'b0001110000000000;
                5'd22: pixel_row = 16'b0011100000000000;
                5'd23: pixel_row = 16'b0011100000000000;
                5'd24: pixel_row = 16'b0111000000000000;
                5'd25: pixel_row = 16'b0111000000000000;
                5'd26: pixel_row = 16'b1110000000000000;
                5'd27: pixel_row = 16'b1110000000000000;
                5'd28: pixel_row = 16'b1110000000000000;
                5'd29: pixel_row = 16'b1100000000000000;
                5'd30: pixel_row = 16'b1100000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '8' - ASCII 56
        //=====================================================
        6'd8: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0011111111111100;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111100000011110;
                5'd4:  pixel_row = 16'b1111000000001111;
                5'd5:  pixel_row = 16'b1110000000000111;
                5'd6:  pixel_row = 16'b1110000000000111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1111000000001111;
                5'd9:  pixel_row = 16'b0111100000011110;
                5'd10: pixel_row = 16'b0011111111111100;
                5'd11: pixel_row = 16'b0001111111111000;
                5'd12: pixel_row = 16'b0011111111111100;
                5'd13: pixel_row = 16'b0111100000011110;
                5'd14: pixel_row = 16'b1111000000001111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                5'd17: pixel_row = 16'b1110000000000111;
                5'd18: pixel_row = 16'b1110000000000111;
                5'd19: pixel_row = 16'b1110000000000111;
                5'd20: pixel_row = 16'b1110000000000111;
                5'd21: pixel_row = 16'b1110000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1111000000001111;
                5'd24: pixel_row = 16'b0111100000011110;
                5'd25: pixel_row = 16'b0111110000111110;
                5'd26: pixel_row = 16'b0011111111111100;
                5'd27: pixel_row = 16'b0001111111111000;
                5'd28: pixel_row = 16'b0000111111110000;
                5'd29: pixel_row = 16'b0000011111100000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '9' - ASCII 57
        //=====================================================
        6'd9: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0011111111111100;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111110000111110;
                5'd4:  pixel_row = 16'b1111100000011111;
                5'd5:  pixel_row = 16'b1111000000001111;
                5'd6:  pixel_row = 16'b1110000000000111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1110000000000111;
                5'd9:  pixel_row = 16'b1110000000000111;
                5'd10: pixel_row = 16'b1110000000000111;
                5'd11: pixel_row = 16'b1110000000000111;
                5'd12: pixel_row = 16'b1110000000000111;
                5'd13: pixel_row = 16'b1111000000000111;
                5'd14: pixel_row = 16'b1111100000001111;
                5'd15: pixel_row = 16'b0111110000011111;
                5'd16: pixel_row = 16'b0111111111111111;
                5'd17: pixel_row = 16'b0011111111110111;
                5'd18: pixel_row = 16'b0001111110000111;
                5'd19: pixel_row = 16'b0000000000000111;
                5'd20: pixel_row = 16'b0000000000000111;
                5'd21: pixel_row = 16'b0000000000001111;
                5'd22: pixel_row = 16'b0000000000001110;
                5'd23: pixel_row = 16'b0000000000011110;
                5'd24: pixel_row = 16'b0000000000111100;
                5'd25: pixel_row = 16'b0000000001111000;
                5'd26: pixel_row = 16'b0111110011110000;
                5'd27: pixel_row = 16'b0111111111100000;
                5'd28: pixel_row = 16'b0011111111000000;
                5'd29: pixel_row = 16'b0001111110000000;
                5'd30: pixel_row = 16'b0000111100000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '.' - 点号 (ASCII 46)
        //=====================================================
        6'd10: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000000000000000;
                5'd5:  pixel_row = 16'b0000000000000000;
                5'd6:  pixel_row = 16'b0000000000000000;
                5'd7:  pixel_row = 16'b0000000000000000;
                5'd8:  pixel_row = 16'b0000000000000000;
                5'd9:  pixel_row = 16'b0000000000000000;
                5'd10: pixel_row = 16'b0000000000000000;
                5'd11: pixel_row = 16'b0000000000000000;
                5'd12: pixel_row = 16'b0000000000000000;
                5'd13: pixel_row = 16'b0000000000000000;
                5'd14: pixel_row = 16'b0000000000000000;
                5'd15: pixel_row = 16'b0000000000000000;
                5'd16: pixel_row = 16'b0000000000000000;
                5'd17: pixel_row = 16'b0000000000000000;
                5'd18: pixel_row = 16'b0000000000000000;
                5'd19: pixel_row = 16'b0000000000000000;
                5'd20: pixel_row = 16'b0000000000000000;
                5'd21: pixel_row = 16'b0000000000000000;
                5'd22: pixel_row = 16'b0000000000000000;
                5'd23: pixel_row = 16'b0000000000000000;
                5'd24: pixel_row = 16'b0000011111000000;
                5'd25: pixel_row = 16'b0000011111000000;
                5'd26: pixel_row = 16'b0000011111000000;
                5'd27: pixel_row = 16'b0000011111000000;
                5'd28: pixel_row = 16'b0000011111000000;
                5'd29: pixel_row = 16'b0000011111000000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // ':' - 冒号 (ASCII 58)
        //=====================================================
        6'd11: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000000000000000;
                5'd5:  pixel_row = 16'b0000000000000000;
                5'd6:  pixel_row = 16'b0000000000000000;
                5'd7:  pixel_row = 16'b0000011111000000;
                5'd8:  pixel_row = 16'b0000011111000000;
                5'd9:  pixel_row = 16'b0000011111000000;
                5'd10: pixel_row = 16'b0000011111000000;
                5'd11: pixel_row = 16'b0000011111000000;
                5'd12: pixel_row = 16'b0000011111000000;
                5'd13: pixel_row = 16'b0000000000000000;
                5'd14: pixel_row = 16'b0000000000000000;
                5'd15: pixel_row = 16'b0000000000000000;
                5'd16: pixel_row = 16'b0000000000000000;
                5'd17: pixel_row = 16'b0000000000000000;
                5'd18: pixel_row = 16'b0000000000000000;
                5'd19: pixel_row = 16'b0000011111000000;
                5'd20: pixel_row = 16'b0000011111000000;
                5'd21: pixel_row = 16'b0000011111000000;
                5'd22: pixel_row = 16'b0000011111000000;
                5'd23: pixel_row = 16'b0000011111000000;
                5'd24: pixel_row = 16'b0000011111000000;
                5'd25: pixel_row = 16'b0000000000000000;
                5'd26: pixel_row = 16'b0000000000000000;
                5'd27: pixel_row = 16'b0000000000000000;
                5'd28: pixel_row = 16'b0000000000000000;
                5'd29: pixel_row = 16'b0000000000000000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '%' - 百分号 (ASCII 37)
        //=====================================================
        6'd12: begin
            case (row)
                5'd0:  pixel_row = 16'b0111000000000110;
                5'd1:  pixel_row = 16'b1101100000001110;
                5'd2:  pixel_row = 16'b1101100000011100;
                5'd3:  pixel_row = 16'b1101100000111000;
                5'd4:  pixel_row = 16'b1101100000110000;
                5'd5:  pixel_row = 16'b0111000001110000;
                5'd6:  pixel_row = 16'b0000000011100000;
                5'd7:  pixel_row = 16'b0000000111000000;
                5'd8:  pixel_row = 16'b0000000110000000;
                5'd9:  pixel_row = 16'b0000001110000000;
                5'd10: pixel_row = 16'b0000011100000000;
                5'd11: pixel_row = 16'b0000011000000000;
                5'd12: pixel_row = 16'b0000111000000000;
                5'd13: pixel_row = 16'b0000110000000000;
                5'd14: pixel_row = 16'b0001110000000000;
                5'd15: pixel_row = 16'b0011100000000000;
                5'd16: pixel_row = 16'b0011000000000000;
                5'd17: pixel_row = 16'b0111000000000000;
                5'd18: pixel_row = 16'b0110000000111000;
                5'd19: pixel_row = 16'b1110000001101100;
                5'd20: pixel_row = 16'b1100000001101100;
                5'd21: pixel_row = 16'b1100000001101100;
                5'd22: pixel_row = 16'b0000000001101100;
                5'd23: pixel_row = 16'b0000000000111000;
                5'd24: pixel_row = 16'b0000000000000000;
                5'd25: pixel_row = 16'b0000000000000000;
                5'd26: pixel_row = 16'b0000000000000000;
                5'd27: pixel_row = 16'b0000000000000000;
                5'd28: pixel_row = 16'b0000000000000000;
                5'd29: pixel_row = 16'b0000000000000000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'H' - 字母H (ASCII 72)
        //=====================================================
        6'd13: begin
            case (row)
                5'd0:  pixel_row = 16'b1110000000000111;
                5'd1:  pixel_row = 16'b1110000000000111;
                5'd2:  pixel_row = 16'b1110000000000111;
                5'd3:  pixel_row = 16'b1110000000000111;
                5'd4:  pixel_row = 16'b1110000000000111;
                5'd5:  pixel_row = 16'b1110000000000111;
                5'd6:  pixel_row = 16'b1110000000000111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1110000000000111;
                5'd9:  pixel_row = 16'b1110000000000111;
                5'd10: pixel_row = 16'b1110000000000111;
                5'd11: pixel_row = 16'b1111111111111111;
                5'd12: pixel_row = 16'b1111111111111111;
                5'd13: pixel_row = 16'b1111111111111111;
                5'd14: pixel_row = 16'b1111111111111111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                5'd17: pixel_row = 16'b1110000000000111;
                5'd18: pixel_row = 16'b1110000000000111;
                5'd19: pixel_row = 16'b1110000000000111;
                5'd20: pixel_row = 16'b1110000000000111;
                5'd21: pixel_row = 16'b1110000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1110000000000111;
                5'd24: pixel_row = 16'b1110000000000111;
                5'd25: pixel_row = 16'b1110000000000111;
                5'd26: pixel_row = 16'b1110000000000111;
                5'd27: pixel_row = 16'b1110000000000111;
                5'd28: pixel_row = 16'b1110000000000111;
                5'd29: pixel_row = 16'b1110000000000111;
                5'd30: pixel_row = 16'b1110000000000111;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'z' - 字母z (ASCII 122)
        //=====================================================
        6'd14: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000000000000000;
                5'd5:  pixel_row = 16'b0111111111111110;
                5'd6:  pixel_row = 16'b0111111111111110;
                5'd7:  pixel_row = 16'b0111111111111110;
                5'd8:  pixel_row = 16'b0000000000111110;
                5'd9:  pixel_row = 16'b0000000001111100;
                5'd10: pixel_row = 16'b0000000011111000;
                5'd11: pixel_row = 16'b0000000111110000;
                5'd12: pixel_row = 16'b0000001111100000;
                5'd13: pixel_row = 16'b0000011111000000;
                5'd14: pixel_row = 16'b0000111110000000;
                5'd15: pixel_row = 16'b0001111100000000;
                5'd16: pixel_row = 16'b0011111000000000;
                5'd17: pixel_row = 16'b0111110000000000;
                5'd18: pixel_row = 16'b0111100000000000;
                5'd19: pixel_row = 16'b1111000000000000;
                5'd20: pixel_row = 16'b1110000000000000;
                5'd21: pixel_row = 16'b1111111111111110;
                5'd22: pixel_row = 16'b1111111111111110;
                5'd23: pixel_row = 16'b1111111111111110;
                5'd24: pixel_row = 16'b0000000000000000;
                5'd25: pixel_row = 16'b0000000000000000;
                5'd26: pixel_row = 16'b0000000000000000;
                5'd27: pixel_row = 16'b0000000000000000;
                5'd28: pixel_row = 16'b0000000000000000;
                5'd29: pixel_row = 16'b0000000000000000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 空格 (ASCII 32)
        //=====================================================
        default: pixel_row = 16'b0000000000000000;
    endcase
end

endmodule
