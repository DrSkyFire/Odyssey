//=============================================================================
// 文件名: ascii_rom_16x32_full.v
// 功能: 完整ASCII字符ROM (16×32像素)
// 字符范围: ASCII 32-126 (空格到~,共95个字符)
// 自动生成: generate_ascii_font.py
// 生成时间: 2025-10-26 22:28:27
//=============================================================================

module ascii_rom_16x32_full (
    input        clk,
    input  [7:0] char_code,   // ASCII码 (32-126有效)
    input  [4:0] char_row,    // 字符行号 (0-31)
    output [15:0] char_data   // 16位字符行数据
);

//=============================================================================
// ROM存储器: 95个字符 × 32行 = 3040行数据
//=============================================================================
reg [15:0] rom [0:3039];

initial begin

    // ASCII 32 (0): ' '
    rom[   0] = 16'b0000000000000000;
    rom[   1] = 16'b0000000000000000;
    rom[   2] = 16'b0000000000000000;
    rom[   3] = 16'b0000000000000000;
    rom[   4] = 16'b0000000000000000;
    rom[   5] = 16'b0000000000000000;
    rom[   6] = 16'b0000000000000000;
    rom[   7] = 16'b0000000000000000;
    rom[   8] = 16'b0000000000000000;
    rom[   9] = 16'b0000000000000000;
    rom[  10] = 16'b0000000000000000;
    rom[  11] = 16'b0000000000000000;
    rom[  12] = 16'b0000000000000000;
    rom[  13] = 16'b0000000000000000;
    rom[  14] = 16'b0000000000000000;
    rom[  15] = 16'b0000000000000000;
    rom[  16] = 16'b0000000000000000;
    rom[  17] = 16'b0000000000000000;
    rom[  18] = 16'b0000000000000000;
    rom[  19] = 16'b0000000000000000;
    rom[  20] = 16'b0000000000000000;
    rom[  21] = 16'b0000000000000000;
    rom[  22] = 16'b0000000000000000;
    rom[  23] = 16'b0000000000000000;
    rom[  24] = 16'b0000000000000000;
    rom[  25] = 16'b0000000000000000;
    rom[  26] = 16'b0000000000000000;
    rom[  27] = 16'b0000000000000000;
    rom[  28] = 16'b0000000000000000;
    rom[  29] = 16'b0000000000000000;
    rom[  30] = 16'b0000000000000000;
    rom[  31] = 16'b0000000000000000;

    // ASCII 33 (1): '!'
    rom[  32] = 16'b0000000000000000;
    rom[  33] = 16'b0000000000000000;
    rom[  34] = 16'b0000000000000000;
    rom[  35] = 16'b0000000000000000;
    rom[  36] = 16'b0000000000000000;
    rom[  37] = 16'b0000000000000000;
    rom[  38] = 16'b0000001100000000;
    rom[  39] = 16'b0000001100000000;
    rom[  40] = 16'b0000001100000000;
    rom[  41] = 16'b0000001100000000;
    rom[  42] = 16'b0000001100000000;
    rom[  43] = 16'b0000001100000000;
    rom[  44] = 16'b0000001100000000;
    rom[  45] = 16'b0000001100000000;
    rom[  46] = 16'b0000001100000000;
    rom[  47] = 16'b0000001100000000;
    rom[  48] = 16'b0000001100000000;
    rom[  49] = 16'b0000001100000000;
    rom[  50] = 16'b0000000000000000;
    rom[  51] = 16'b0000000000000000;
    rom[  52] = 16'b0000001110000000;
    rom[  53] = 16'b0000001110000000;
    rom[  54] = 16'b0000001110000000;
    rom[  55] = 16'b0000000000000000;
    rom[  56] = 16'b0000000000000000;
    rom[  57] = 16'b0000000000000000;
    rom[  58] = 16'b0000000000000000;
    rom[  59] = 16'b0000000000000000;
    rom[  60] = 16'b0000000000000000;
    rom[  61] = 16'b0000000000000000;
    rom[  62] = 16'b0000000000000000;
    rom[  63] = 16'b0000000000000000;

    // ASCII 34 (2): '"'
    rom[  64] = 16'b0000000000000000;
    rom[  65] = 16'b0000000000000000;
    rom[  66] = 16'b0000000000000000;
    rom[  67] = 16'b0000000000000000;
    rom[  68] = 16'b0000000000000000;
    rom[  69] = 16'b0000000000000000;
    rom[  70] = 16'b0000111001110000;
    rom[  71] = 16'b0000111001110000;
    rom[  72] = 16'b0000111001110000;
    rom[  73] = 16'b0000111001110000;
    rom[  74] = 16'b0000111001110000;
    rom[  75] = 16'b0000111001110000;
    rom[  76] = 16'b0000000000000000;
    rom[  77] = 16'b0000000000000000;
    rom[  78] = 16'b0000000000000000;
    rom[  79] = 16'b0000000000000000;
    rom[  80] = 16'b0000000000000000;
    rom[  81] = 16'b0000000000000000;
    rom[  82] = 16'b0000000000000000;
    rom[  83] = 16'b0000000000000000;
    rom[  84] = 16'b0000000000000000;
    rom[  85] = 16'b0000000000000000;
    rom[  86] = 16'b0000000000000000;
    rom[  87] = 16'b0000000000000000;
    rom[  88] = 16'b0000000000000000;
    rom[  89] = 16'b0000000000000000;
    rom[  90] = 16'b0000000000000000;
    rom[  91] = 16'b0000000000000000;
    rom[  92] = 16'b0000000000000000;
    rom[  93] = 16'b0000000000000000;
    rom[  94] = 16'b0000000000000000;
    rom[  95] = 16'b0000000000000000;

    // ASCII 35 (3): '#'
    rom[  96] = 16'b0000000000000000;
    rom[  97] = 16'b0000000000000000;
    rom[  98] = 16'b0000000000000000;
    rom[  99] = 16'b0000000000000000;
    rom[ 100] = 16'b0000000000000000;
    rom[ 101] = 16'b0000000000000000;
    rom[ 102] = 16'b0000000000000000;
    rom[ 103] = 16'b0000000000000000;
    rom[ 104] = 16'b0000000000000000;
    rom[ 105] = 16'b0000001100110000;
    rom[ 106] = 16'b0000001100110000;
    rom[ 107] = 16'b0000001100110000;
    rom[ 108] = 16'b0000001100110000;
    rom[ 109] = 16'b0001111111111100;
    rom[ 110] = 16'b0001111111111100;
    rom[ 111] = 16'b0000011001100000;
    rom[ 112] = 16'b0000011001100000;
    rom[ 113] = 16'b0000011001100000;
    rom[ 114] = 16'b0011111111111000;
    rom[ 115] = 16'b0011111111111000;
    rom[ 116] = 16'b0000111011100000;
    rom[ 117] = 16'b0000110011000000;
    rom[ 118] = 16'b0000110011000000;
    rom[ 119] = 16'b0000110011000000;
    rom[ 120] = 16'b0000000000000000;
    rom[ 121] = 16'b0000000000000000;
    rom[ 122] = 16'b0000000000000000;
    rom[ 123] = 16'b0000000000000000;
    rom[ 124] = 16'b0000000000000000;
    rom[ 125] = 16'b0000000000000000;
    rom[ 126] = 16'b0000000000000000;
    rom[ 127] = 16'b0000000000000000;

    // ASCII 36 (4): '$'
    rom[ 128] = 16'b0000000000000000;
    rom[ 129] = 16'b0000000000000000;
    rom[ 130] = 16'b0000000000000000;
    rom[ 131] = 16'b0000000110000000;
    rom[ 132] = 16'b0000000110000000;
    rom[ 133] = 16'b0000011111100000;
    rom[ 134] = 16'b0001111111100000;
    rom[ 135] = 16'b0011100110000000;
    rom[ 136] = 16'b0011000100000000;
    rom[ 137] = 16'b0011000100000000;
    rom[ 138] = 16'b0011101100000000;
    rom[ 139] = 16'b0001111100000000;
    rom[ 140] = 16'b0000111110000000;
    rom[ 141] = 16'b0000001111000000;
    rom[ 142] = 16'b0000001111100000;
    rom[ 143] = 16'b0000001100110000;
    rom[ 144] = 16'b0000001000110000;
    rom[ 145] = 16'b0000001000110000;
    rom[ 146] = 16'b0010011001110000;
    rom[ 147] = 16'b0011111111100000;
    rom[ 148] = 16'b0001111110000000;
    rom[ 149] = 16'b0000011000000000;
    rom[ 150] = 16'b0000011000000000;
    rom[ 151] = 16'b0000011000000000;
    rom[ 152] = 16'b0000000000000000;
    rom[ 153] = 16'b0000000000000000;
    rom[ 154] = 16'b0000000000000000;
    rom[ 155] = 16'b0000000000000000;
    rom[ 156] = 16'b0000000000000000;
    rom[ 157] = 16'b0000000000000000;
    rom[ 158] = 16'b0000000000000000;
    rom[ 159] = 16'b0000000000000000;

    // ASCII 37 (5): '%'
    rom[ 160] = 16'b0000000000000000;
    rom[ 161] = 16'b0000000000000000;
    rom[ 162] = 16'b0000000000000000;
    rom[ 163] = 16'b0000000000000000;
    rom[ 164] = 16'b0000000000000000;
    rom[ 165] = 16'b0000000000000000;
    rom[ 166] = 16'b0001111000001100;
    rom[ 167] = 16'b0011111100011000;
    rom[ 168] = 16'b0110001100110000;
    rom[ 169] = 16'b0110001100110000;
    rom[ 170] = 16'b0110001101100000;
    rom[ 171] = 16'b0111111011000000;
    rom[ 172] = 16'b0011110011000000;
    rom[ 173] = 16'b0000000110000000;
    rom[ 174] = 16'b0000001100000000;
    rom[ 175] = 16'b0000001100000000;
    rom[ 176] = 16'b0000011001111000;
    rom[ 177] = 16'b0000011011111100;
    rom[ 178] = 16'b0000110110001100;
    rom[ 179] = 16'b0001100110001100;
    rom[ 180] = 16'b0001100110001100;
    rom[ 181] = 16'b0011000111111000;
    rom[ 182] = 16'b0110000011110000;
    rom[ 183] = 16'b0000000000000000;
    rom[ 184] = 16'b0000000000000000;
    rom[ 185] = 16'b0000000000000000;
    rom[ 186] = 16'b0000000000000000;
    rom[ 187] = 16'b0000000000000000;
    rom[ 188] = 16'b0000000000000000;
    rom[ 189] = 16'b0000000000000000;
    rom[ 190] = 16'b0000000000000000;
    rom[ 191] = 16'b0000000000000000;

    // ASCII 38 (6): '&'
    rom[ 192] = 16'b0000000000000000;
    rom[ 193] = 16'b0000000000000000;
    rom[ 194] = 16'b0000000000000000;
    rom[ 195] = 16'b0000000000000000;
    rom[ 196] = 16'b0000000000000000;
    rom[ 197] = 16'b0000000000000000;
    rom[ 198] = 16'b0000011110000000;
    rom[ 199] = 16'b0000111111000000;
    rom[ 200] = 16'b0001110011100000;
    rom[ 201] = 16'b0001100001100000;
    rom[ 202] = 16'b0001100001100000;
    rom[ 203] = 16'b0001100011100000;
    rom[ 204] = 16'b0001110111000000;
    rom[ 205] = 16'b0000111110000000;
    rom[ 206] = 16'b0000111100000000;
    rom[ 207] = 16'b0001111100011000;
    rom[ 208] = 16'b0011101110011000;
    rom[ 209] = 16'b0011000111011000;
    rom[ 210] = 16'b0011000011110000;
    rom[ 211] = 16'b0011000001110000;
    rom[ 212] = 16'b0011100011110000;
    rom[ 213] = 16'b0001111111111000;
    rom[ 214] = 16'b0000111110011100;
    rom[ 215] = 16'b0000000000000000;
    rom[ 216] = 16'b0000000000000000;
    rom[ 217] = 16'b0000000000000000;
    rom[ 218] = 16'b0000000000000000;
    rom[ 219] = 16'b0000000000000000;
    rom[ 220] = 16'b0000000000000000;
    rom[ 221] = 16'b0000000000000000;
    rom[ 222] = 16'b0000000000000000;
    rom[ 223] = 16'b0000000000000000;

    // ASCII 39 (7): "'"
    rom[ 224] = 16'b0000000000000000;
    rom[ 225] = 16'b0000000000000000;
    rom[ 226] = 16'b0000000000000000;
    rom[ 227] = 16'b0000000000000000;
    rom[ 228] = 16'b0000000000000000;
    rom[ 229] = 16'b0000000000000000;
    rom[ 230] = 16'b0000001110000000;
    rom[ 231] = 16'b0000001110000000;
    rom[ 232] = 16'b0000001110000000;
    rom[ 233] = 16'b0000001110000000;
    rom[ 234] = 16'b0000001110000000;
    rom[ 235] = 16'b0000001110000000;
    rom[ 236] = 16'b0000000000000000;
    rom[ 237] = 16'b0000000000000000;
    rom[ 238] = 16'b0000000000000000;
    rom[ 239] = 16'b0000000000000000;
    rom[ 240] = 16'b0000000000000000;
    rom[ 241] = 16'b0000000000000000;
    rom[ 242] = 16'b0000000000000000;
    rom[ 243] = 16'b0000000000000000;
    rom[ 244] = 16'b0000000000000000;
    rom[ 245] = 16'b0000000000000000;
    rom[ 246] = 16'b0000000000000000;
    rom[ 247] = 16'b0000000000000000;
    rom[ 248] = 16'b0000000000000000;
    rom[ 249] = 16'b0000000000000000;
    rom[ 250] = 16'b0000000000000000;
    rom[ 251] = 16'b0000000000000000;
    rom[ 252] = 16'b0000000000000000;
    rom[ 253] = 16'b0000000000000000;
    rom[ 254] = 16'b0000000000000000;
    rom[ 255] = 16'b0000000000000000;

    // ASCII 40 (8): '('
    rom[ 256] = 16'b0000000000000000;
    rom[ 257] = 16'b0000000000000000;
    rom[ 258] = 16'b0000000000000000;
    rom[ 259] = 16'b0000000000000000;
    rom[ 260] = 16'b0000000000100000;
    rom[ 261] = 16'b0000000001110000;
    rom[ 262] = 16'b0000000011100000;
    rom[ 263] = 16'b0000000111000000;
    rom[ 264] = 16'b0000000110000000;
    rom[ 265] = 16'b0000001100000000;
    rom[ 266] = 16'b0000001100000000;
    rom[ 267] = 16'b0000001100000000;
    rom[ 268] = 16'b0000011000000000;
    rom[ 269] = 16'b0000011000000000;
    rom[ 270] = 16'b0000011000000000;
    rom[ 271] = 16'b0000011000000000;
    rom[ 272] = 16'b0000011000000000;
    rom[ 273] = 16'b0000011000000000;
    rom[ 274] = 16'b0000011100000000;
    rom[ 275] = 16'b0000001100000000;
    rom[ 276] = 16'b0000001100000000;
    rom[ 277] = 16'b0000000110000000;
    rom[ 278] = 16'b0000000111000000;
    rom[ 279] = 16'b0000000011100000;
    rom[ 280] = 16'b0000000001110000;
    rom[ 281] = 16'b0000000000100000;
    rom[ 282] = 16'b0000000000000000;
    rom[ 283] = 16'b0000000000000000;
    rom[ 284] = 16'b0000000000000000;
    rom[ 285] = 16'b0000000000000000;
    rom[ 286] = 16'b0000000000000000;
    rom[ 287] = 16'b0000000000000000;

    // ASCII 41 (9): ')'
    rom[ 288] = 16'b0000000000000000;
    rom[ 289] = 16'b0000000000000000;
    rom[ 290] = 16'b0000000000000000;
    rom[ 291] = 16'b0000000000000000;
    rom[ 292] = 16'b0000010000000000;
    rom[ 293] = 16'b0000111000000000;
    rom[ 294] = 16'b0000011100000000;
    rom[ 295] = 16'b0000001110000000;
    rom[ 296] = 16'b0000000110000000;
    rom[ 297] = 16'b0000000011000000;
    rom[ 298] = 16'b0000000011000000;
    rom[ 299] = 16'b0000000011100000;
    rom[ 300] = 16'b0000000001100000;
    rom[ 301] = 16'b0000000001100000;
    rom[ 302] = 16'b0000000001100000;
    rom[ 303] = 16'b0000000001100000;
    rom[ 304] = 16'b0000000001100000;
    rom[ 305] = 16'b0000000001100000;
    rom[ 306] = 16'b0000000011000000;
    rom[ 307] = 16'b0000000011000000;
    rom[ 308] = 16'b0000000011000000;
    rom[ 309] = 16'b0000000110000000;
    rom[ 310] = 16'b0000001110000000;
    rom[ 311] = 16'b0000011100000000;
    rom[ 312] = 16'b0000111000000000;
    rom[ 313] = 16'b0000010000000000;
    rom[ 314] = 16'b0000000000000000;
    rom[ 315] = 16'b0000000000000000;
    rom[ 316] = 16'b0000000000000000;
    rom[ 317] = 16'b0000000000000000;
    rom[ 318] = 16'b0000000000000000;
    rom[ 319] = 16'b0000000000000000;

    // ASCII 42 (10): '*'
    rom[ 320] = 16'b0000000000000000;
    rom[ 321] = 16'b0000000000000000;
    rom[ 322] = 16'b0000000000000000;
    rom[ 323] = 16'b0000000000000000;
    rom[ 324] = 16'b0000000000000000;
    rom[ 325] = 16'b0000000000000000;
    rom[ 326] = 16'b0000000110000000;
    rom[ 327] = 16'b0000000110000000;
    rom[ 328] = 16'b0000100110010000;
    rom[ 329] = 16'b0001110110111000;
    rom[ 330] = 16'b0000001111000000;
    rom[ 331] = 16'b0000001111000000;
    rom[ 332] = 16'b0001110110111000;
    rom[ 333] = 16'b0001100110011000;
    rom[ 334] = 16'b0000000110000000;
    rom[ 335] = 16'b0000000110000000;
    rom[ 336] = 16'b0000000000000000;
    rom[ 337] = 16'b0000000000000000;
    rom[ 338] = 16'b0000000000000000;
    rom[ 339] = 16'b0000000000000000;
    rom[ 340] = 16'b0000000000000000;
    rom[ 341] = 16'b0000000000000000;
    rom[ 342] = 16'b0000000000000000;
    rom[ 343] = 16'b0000000000000000;
    rom[ 344] = 16'b0000000000000000;
    rom[ 345] = 16'b0000000000000000;
    rom[ 346] = 16'b0000000000000000;
    rom[ 347] = 16'b0000000000000000;
    rom[ 348] = 16'b0000000000000000;
    rom[ 349] = 16'b0000000000000000;
    rom[ 350] = 16'b0000000000000000;
    rom[ 351] = 16'b0000000000000000;

    // ASCII 43 (11): '+'
    rom[ 352] = 16'b0000000000000000;
    rom[ 353] = 16'b0000000000000000;
    rom[ 354] = 16'b0000000000000000;
    rom[ 355] = 16'b0000000000000000;
    rom[ 356] = 16'b0000000000000000;
    rom[ 357] = 16'b0000000000000000;
    rom[ 358] = 16'b0000000000000000;
    rom[ 359] = 16'b0000000000000000;
    rom[ 360] = 16'b0000000000000000;
    rom[ 361] = 16'b0000000000000000;
    rom[ 362] = 16'b0000000000000000;
    rom[ 363] = 16'b0000000000000000;
    rom[ 364] = 16'b0000000110000000;
    rom[ 365] = 16'b0000000110000000;
    rom[ 366] = 16'b0000000110000000;
    rom[ 367] = 16'b0000000110000000;
    rom[ 368] = 16'b0000000110000000;
    rom[ 369] = 16'b0011111111111100;
    rom[ 370] = 16'b0011111111111100;
    rom[ 371] = 16'b0000000110000000;
    rom[ 372] = 16'b0000000110000000;
    rom[ 373] = 16'b0000000110000000;
    rom[ 374] = 16'b0000000110000000;
    rom[ 375] = 16'b0000000110000000;
    rom[ 376] = 16'b0000000000000000;
    rom[ 377] = 16'b0000000000000000;
    rom[ 378] = 16'b0000000000000000;
    rom[ 379] = 16'b0000000000000000;
    rom[ 380] = 16'b0000000000000000;
    rom[ 381] = 16'b0000000000000000;
    rom[ 382] = 16'b0000000000000000;
    rom[ 383] = 16'b0000000000000000;

    // ASCII 44 (12): ','
    rom[ 384] = 16'b0000000000000000;
    rom[ 385] = 16'b0000000000000000;
    rom[ 386] = 16'b0000000000000000;
    rom[ 387] = 16'b0000000000000000;
    rom[ 388] = 16'b0000000000000000;
    rom[ 389] = 16'b0000000000000000;
    rom[ 390] = 16'b0000000000000000;
    rom[ 391] = 16'b0000000000000000;
    rom[ 392] = 16'b0000000000000000;
    rom[ 393] = 16'b0000000000000000;
    rom[ 394] = 16'b0000000000000000;
    rom[ 395] = 16'b0000000000000000;
    rom[ 396] = 16'b0000000000000000;
    rom[ 397] = 16'b0000000000000000;
    rom[ 398] = 16'b0000000000000000;
    rom[ 399] = 16'b0000000000000000;
    rom[ 400] = 16'b0000000000000000;
    rom[ 401] = 16'b0000000000000000;
    rom[ 402] = 16'b0000000000000000;
    rom[ 403] = 16'b0000000000000000;
    rom[ 404] = 16'b0000000000000000;
    rom[ 405] = 16'b0000000000000000;
    rom[ 406] = 16'b0000000000000000;
    rom[ 407] = 16'b0000000000000000;
    rom[ 408] = 16'b0000001110000000;
    rom[ 409] = 16'b0000001111000000;
    rom[ 410] = 16'b0000001111000000;
    rom[ 411] = 16'b0000000111000000;
    rom[ 412] = 16'b0000000111000000;
    rom[ 413] = 16'b0000001110000000;
    rom[ 414] = 16'b0000111100000000;
    rom[ 415] = 16'b0000111000000000;

    // ASCII 45 (13): '-'
    rom[ 416] = 16'b0000000000000000;
    rom[ 417] = 16'b0000000000000000;
    rom[ 418] = 16'b0000000000000000;
    rom[ 419] = 16'b0000000000000000;
    rom[ 420] = 16'b0000000000000000;
    rom[ 421] = 16'b0000000000000000;
    rom[ 422] = 16'b0000000000000000;
    rom[ 423] = 16'b0000000000000000;
    rom[ 424] = 16'b0000000000000000;
    rom[ 425] = 16'b0000000000000000;
    rom[ 426] = 16'b0000000000000000;
    rom[ 427] = 16'b0000000000000000;
    rom[ 428] = 16'b0000000000000000;
    rom[ 429] = 16'b0000000000000000;
    rom[ 430] = 16'b0000000000000000;
    rom[ 431] = 16'b0000000000000000;
    rom[ 432] = 16'b0000000000000000;
    rom[ 433] = 16'b0000000000000000;
    rom[ 434] = 16'b0000000000000000;
    rom[ 435] = 16'b0000000000000000;
    rom[ 436] = 16'b0000000000000000;
    rom[ 437] = 16'b0000111111100000;
    rom[ 438] = 16'b0000111111100000;
    rom[ 439] = 16'b0000000000000000;
    rom[ 440] = 16'b0000000000000000;
    rom[ 441] = 16'b0000000000000000;
    rom[ 442] = 16'b0000000000000000;
    rom[ 443] = 16'b0000000000000000;
    rom[ 444] = 16'b0000000000000000;
    rom[ 445] = 16'b0000000000000000;
    rom[ 446] = 16'b0000000000000000;
    rom[ 447] = 16'b0000000000000000;

    // ASCII 46 (14): '.'
    rom[ 448] = 16'b0000000000000000;
    rom[ 449] = 16'b0000000000000000;
    rom[ 450] = 16'b0000000000000000;
    rom[ 451] = 16'b0000000000000000;
    rom[ 452] = 16'b0000000000000000;
    rom[ 453] = 16'b0000000000000000;
    rom[ 454] = 16'b0000000000000000;
    rom[ 455] = 16'b0000000000000000;
    rom[ 456] = 16'b0000000000000000;
    rom[ 457] = 16'b0000000000000000;
    rom[ 458] = 16'b0000000000000000;
    rom[ 459] = 16'b0000000000000000;
    rom[ 460] = 16'b0000000000000000;
    rom[ 461] = 16'b0000000000000000;
    rom[ 462] = 16'b0000000000000000;
    rom[ 463] = 16'b0000000000000000;
    rom[ 464] = 16'b0000000000000000;
    rom[ 465] = 16'b0000000000000000;
    rom[ 466] = 16'b0000000000000000;
    rom[ 467] = 16'b0000000000000000;
    rom[ 468] = 16'b0000000000000000;
    rom[ 469] = 16'b0000000000000000;
    rom[ 470] = 16'b0000000000000000;
    rom[ 471] = 16'b0000000000000000;
    rom[ 472] = 16'b0000000000000000;
    rom[ 473] = 16'b0000000000000000;
    rom[ 474] = 16'b0000000110000000;
    rom[ 475] = 16'b0000001111000000;
    rom[ 476] = 16'b0000001111000000;
    rom[ 477] = 16'b0000000110000000;
    rom[ 478] = 16'b0000000000000000;
    rom[ 479] = 16'b0000000000000000;

    // ASCII 47 (15): '/'
    rom[ 480] = 16'b0000000000000000;
    rom[ 481] = 16'b0000000000000000;
    rom[ 482] = 16'b0000000000000000;
    rom[ 483] = 16'b0000000000000000;
    rom[ 484] = 16'b0000000000000000;
    rom[ 485] = 16'b0000000000110000;
    rom[ 486] = 16'b0000000001100000;
    rom[ 487] = 16'b0000000001100000;
    rom[ 488] = 16'b0000000001100000;
    rom[ 489] = 16'b0000000011000000;
    rom[ 490] = 16'b0000000011000000;
    rom[ 491] = 16'b0000000110000000;
    rom[ 492] = 16'b0000000110000000;
    rom[ 493] = 16'b0000000110000000;
    rom[ 494] = 16'b0000001100000000;
    rom[ 495] = 16'b0000001100000000;
    rom[ 496] = 16'b0000011000000000;
    rom[ 497] = 16'b0000011000000000;
    rom[ 498] = 16'b0000011000000000;
    rom[ 499] = 16'b0000110000000000;
    rom[ 500] = 16'b0000110000000000;
    rom[ 501] = 16'b0001100000000000;
    rom[ 502] = 16'b0001100000000000;
    rom[ 503] = 16'b0001100000000000;
    rom[ 504] = 16'b0011000000000000;
    rom[ 505] = 16'b0000000000000000;
    rom[ 506] = 16'b0000000000000000;
    rom[ 507] = 16'b0000000000000000;
    rom[ 508] = 16'b0000000000000000;
    rom[ 509] = 16'b0000000000000000;
    rom[ 510] = 16'b0000000000000000;
    rom[ 511] = 16'b0000000000000000;

    // ASCII 48 (16): '0'
    rom[ 512] = 16'b0000000000000000;
    rom[ 513] = 16'b0000000000000000;
    rom[ 514] = 16'b0000000000000000;
    rom[ 515] = 16'b0000000000000000;
    rom[ 516] = 16'b0000000000000000;
    rom[ 517] = 16'b0000000000000000;
    rom[ 518] = 16'b0000000000000000;
    rom[ 519] = 16'b0000000000000000;
    rom[ 520] = 16'b0000000000000000;
    rom[ 521] = 16'b0000011111000000;
    rom[ 522] = 16'b0000111111100000;
    rom[ 523] = 16'b0001110001110000;
    rom[ 524] = 16'b0001100000110000;
    rom[ 525] = 16'b0011000000111000;
    rom[ 526] = 16'b0011000001111000;
    rom[ 527] = 16'b0011000111011000;
    rom[ 528] = 16'b0011001110011000;
    rom[ 529] = 16'b0011011100011000;
    rom[ 530] = 16'b0011110000011000;
    rom[ 531] = 16'b0011100000011000;
    rom[ 532] = 16'b0001100000110000;
    rom[ 533] = 16'b0001110001110000;
    rom[ 534] = 16'b0000111111100000;
    rom[ 535] = 16'b0000011111000000;
    rom[ 536] = 16'b0000000000000000;
    rom[ 537] = 16'b0000000000000000;
    rom[ 538] = 16'b0000000000000000;
    rom[ 539] = 16'b0000000000000000;
    rom[ 540] = 16'b0000000000000000;
    rom[ 541] = 16'b0000000000000000;
    rom[ 542] = 16'b0000000000000000;
    rom[ 543] = 16'b0000000000000000;

    // ASCII 49 (17): '1'
    rom[ 544] = 16'b0000000000000000;
    rom[ 545] = 16'b0000000000000000;
    rom[ 546] = 16'b0000000000000000;
    rom[ 547] = 16'b0000000000000000;
    rom[ 548] = 16'b0000000000000000;
    rom[ 549] = 16'b0000000000000000;
    rom[ 550] = 16'b0000000000000000;
    rom[ 551] = 16'b0000000000000000;
    rom[ 552] = 16'b0000000000000000;
    rom[ 553] = 16'b0000001110000000;
    rom[ 554] = 16'b0000111110000000;
    rom[ 555] = 16'b0001110110000000;
    rom[ 556] = 16'b0001100110000000;
    rom[ 557] = 16'b0000000110000000;
    rom[ 558] = 16'b0000000110000000;
    rom[ 559] = 16'b0000000110000000;
    rom[ 560] = 16'b0000000110000000;
    rom[ 561] = 16'b0000000110000000;
    rom[ 562] = 16'b0000000110000000;
    rom[ 563] = 16'b0000000110000000;
    rom[ 564] = 16'b0000000110000000;
    rom[ 565] = 16'b0000000110000000;
    rom[ 566] = 16'b0001111111111000;
    rom[ 567] = 16'b0001111111111000;
    rom[ 568] = 16'b0000000000000000;
    rom[ 569] = 16'b0000000000000000;
    rom[ 570] = 16'b0000000000000000;
    rom[ 571] = 16'b0000000000000000;
    rom[ 572] = 16'b0000000000000000;
    rom[ 573] = 16'b0000000000000000;
    rom[ 574] = 16'b0000000000000000;
    rom[ 575] = 16'b0000000000000000;

    // ASCII 50 (18): '2'
    rom[ 576] = 16'b0000000000000000;
    rom[ 577] = 16'b0000000000000000;
    rom[ 578] = 16'b0000000000000000;
    rom[ 579] = 16'b0000000000000000;
    rom[ 580] = 16'b0000000000000000;
    rom[ 581] = 16'b0000000000000000;
    rom[ 582] = 16'b0000000000000000;
    rom[ 583] = 16'b0000000000000000;
    rom[ 584] = 16'b0000000000000000;
    rom[ 585] = 16'b0000011111000000;
    rom[ 586] = 16'b0000111111100000;
    rom[ 587] = 16'b0001110001110000;
    rom[ 588] = 16'b0000100000110000;
    rom[ 589] = 16'b0000000000110000;
    rom[ 590] = 16'b0000000000110000;
    rom[ 591] = 16'b0000000001110000;
    rom[ 592] = 16'b0000000001100000;
    rom[ 593] = 16'b0000000011000000;
    rom[ 594] = 16'b0000000110000000;
    rom[ 595] = 16'b0000001100000000;
    rom[ 596] = 16'b0000011000000000;
    rom[ 597] = 16'b0000111000000000;
    rom[ 598] = 16'b0001111111111000;
    rom[ 599] = 16'b0001111111111000;
    rom[ 600] = 16'b0000000000000000;
    rom[ 601] = 16'b0000000000000000;
    rom[ 602] = 16'b0000000000000000;
    rom[ 603] = 16'b0000000000000000;
    rom[ 604] = 16'b0000000000000000;
    rom[ 605] = 16'b0000000000000000;
    rom[ 606] = 16'b0000000000000000;
    rom[ 607] = 16'b0000000000000000;

    // ASCII 51 (19): '3'
    rom[ 608] = 16'b0000000000000000;
    rom[ 609] = 16'b0000000000000000;
    rom[ 610] = 16'b0000000000000000;
    rom[ 611] = 16'b0000000000000000;
    rom[ 612] = 16'b0000000000000000;
    rom[ 613] = 16'b0000000000000000;
    rom[ 614] = 16'b0000000000000000;
    rom[ 615] = 16'b0000000000000000;
    rom[ 616] = 16'b0000000000000000;
    rom[ 617] = 16'b0000111110000000;
    rom[ 618] = 16'b0001111111000000;
    rom[ 619] = 16'b0001000011100000;
    rom[ 620] = 16'b0000000001100000;
    rom[ 621] = 16'b0000000001100000;
    rom[ 622] = 16'b0000000011000000;
    rom[ 623] = 16'b0000011110000000;
    rom[ 624] = 16'b0000011111100000;
    rom[ 625] = 16'b0000000001110000;
    rom[ 626] = 16'b0000000000110000;
    rom[ 627] = 16'b0000000000110000;
    rom[ 628] = 16'b0000000000110000;
    rom[ 629] = 16'b0000000001100000;
    rom[ 630] = 16'b0001111111100000;
    rom[ 631] = 16'b0001111110000000;
    rom[ 632] = 16'b0000000000000000;
    rom[ 633] = 16'b0000000000000000;
    rom[ 634] = 16'b0000000000000000;
    rom[ 635] = 16'b0000000000000000;
    rom[ 636] = 16'b0000000000000000;
    rom[ 637] = 16'b0000000000000000;
    rom[ 638] = 16'b0000000000000000;
    rom[ 639] = 16'b0000000000000000;

    // ASCII 52 (20): '4'
    rom[ 640] = 16'b0000000000000000;
    rom[ 641] = 16'b0000000000000000;
    rom[ 642] = 16'b0000000000000000;
    rom[ 643] = 16'b0000000000000000;
    rom[ 644] = 16'b0000000000000000;
    rom[ 645] = 16'b0000000000000000;
    rom[ 646] = 16'b0000000000000000;
    rom[ 647] = 16'b0000000000000000;
    rom[ 648] = 16'b0000000000000000;
    rom[ 649] = 16'b0000000011100000;
    rom[ 650] = 16'b0000000111100000;
    rom[ 651] = 16'b0000000111100000;
    rom[ 652] = 16'b0000001101100000;
    rom[ 653] = 16'b0000011001100000;
    rom[ 654] = 16'b0000011001100000;
    rom[ 655] = 16'b0000110001100000;
    rom[ 656] = 16'b0000110001100000;
    rom[ 657] = 16'b0001100001100000;
    rom[ 658] = 16'b0011000001100000;
    rom[ 659] = 16'b0011111111111100;
    rom[ 660] = 16'b0011111111111100;
    rom[ 661] = 16'b0000000001100000;
    rom[ 662] = 16'b0000000001100000;
    rom[ 663] = 16'b0000000001100000;
    rom[ 664] = 16'b0000000000000000;
    rom[ 665] = 16'b0000000000000000;
    rom[ 666] = 16'b0000000000000000;
    rom[ 667] = 16'b0000000000000000;
    rom[ 668] = 16'b0000000000000000;
    rom[ 669] = 16'b0000000000000000;
    rom[ 670] = 16'b0000000000000000;
    rom[ 671] = 16'b0000000000000000;

    // ASCII 53 (21): '5'
    rom[ 672] = 16'b0000000000000000;
    rom[ 673] = 16'b0000000000000000;
    rom[ 674] = 16'b0000000000000000;
    rom[ 675] = 16'b0000000000000000;
    rom[ 676] = 16'b0000000000000000;
    rom[ 677] = 16'b0000000000000000;
    rom[ 678] = 16'b0000000000000000;
    rom[ 679] = 16'b0000000000000000;
    rom[ 680] = 16'b0000000000000000;
    rom[ 681] = 16'b0001111111100000;
    rom[ 682] = 16'b0001111111100000;
    rom[ 683] = 16'b0001100000000000;
    rom[ 684] = 16'b0001100000000000;
    rom[ 685] = 16'b0001100000000000;
    rom[ 686] = 16'b0001100000000000;
    rom[ 687] = 16'b0001111111000000;
    rom[ 688] = 16'b0001111111100000;
    rom[ 689] = 16'b0000000001110000;
    rom[ 690] = 16'b0000000000110000;
    rom[ 691] = 16'b0000000000110000;
    rom[ 692] = 16'b0000000000110000;
    rom[ 693] = 16'b0000000001100000;
    rom[ 694] = 16'b0001111111000000;
    rom[ 695] = 16'b0001111110000000;
    rom[ 696] = 16'b0000000000000000;
    rom[ 697] = 16'b0000000000000000;
    rom[ 698] = 16'b0000000000000000;
    rom[ 699] = 16'b0000000000000000;
    rom[ 700] = 16'b0000000000000000;
    rom[ 701] = 16'b0000000000000000;
    rom[ 702] = 16'b0000000000000000;
    rom[ 703] = 16'b0000000000000000;

    // ASCII 54 (22): '6'
    rom[ 704] = 16'b0000000000000000;
    rom[ 705] = 16'b0000000000000000;
    rom[ 706] = 16'b0000000000000000;
    rom[ 707] = 16'b0000000000000000;
    rom[ 708] = 16'b0000000000000000;
    rom[ 709] = 16'b0000000000000000;
    rom[ 710] = 16'b0000000000000000;
    rom[ 711] = 16'b0000000000000000;
    rom[ 712] = 16'b0000000000000000;
    rom[ 713] = 16'b0000001111100000;
    rom[ 714] = 16'b0000111111100000;
    rom[ 715] = 16'b0000111000000000;
    rom[ 716] = 16'b0001100000000000;
    rom[ 717] = 16'b0001000000000000;
    rom[ 718] = 16'b0011000000000000;
    rom[ 719] = 16'b0011011111000000;
    rom[ 720] = 16'b0011111111100000;
    rom[ 721] = 16'b0011100001110000;
    rom[ 722] = 16'b0011000000110000;
    rom[ 723] = 16'b0011000000110000;
    rom[ 724] = 16'b0011000000110000;
    rom[ 725] = 16'b0001100001100000;
    rom[ 726] = 16'b0001111111100000;
    rom[ 727] = 16'b0000011110000000;
    rom[ 728] = 16'b0000000000000000;
    rom[ 729] = 16'b0000000000000000;
    rom[ 730] = 16'b0000000000000000;
    rom[ 731] = 16'b0000000000000000;
    rom[ 732] = 16'b0000000000000000;
    rom[ 733] = 16'b0000000000000000;
    rom[ 734] = 16'b0000000000000000;
    rom[ 735] = 16'b0000000000000000;

    // ASCII 55 (23): '7'
    rom[ 736] = 16'b0000000000000000;
    rom[ 737] = 16'b0000000000000000;
    rom[ 738] = 16'b0000000000000000;
    rom[ 739] = 16'b0000000000000000;
    rom[ 740] = 16'b0000000000000000;
    rom[ 741] = 16'b0000000000000000;
    rom[ 742] = 16'b0000000000000000;
    rom[ 743] = 16'b0000000000000000;
    rom[ 744] = 16'b0000000000000000;
    rom[ 745] = 16'b0011111111110000;
    rom[ 746] = 16'b0011111111110000;
    rom[ 747] = 16'b0000000000110000;
    rom[ 748] = 16'b0000000001100000;
    rom[ 749] = 16'b0000000001100000;
    rom[ 750] = 16'b0000000011000000;
    rom[ 751] = 16'b0000000011000000;
    rom[ 752] = 16'b0000000110000000;
    rom[ 753] = 16'b0000000110000000;
    rom[ 754] = 16'b0000001100000000;
    rom[ 755] = 16'b0000001100000000;
    rom[ 756] = 16'b0000011000000000;
    rom[ 757] = 16'b0000011000000000;
    rom[ 758] = 16'b0000111000000000;
    rom[ 759] = 16'b0000110000000000;
    rom[ 760] = 16'b0000000000000000;
    rom[ 761] = 16'b0000000000000000;
    rom[ 762] = 16'b0000000000000000;
    rom[ 763] = 16'b0000000000000000;
    rom[ 764] = 16'b0000000000000000;
    rom[ 765] = 16'b0000000000000000;
    rom[ 766] = 16'b0000000000000000;
    rom[ 767] = 16'b0000000000000000;

    // ASCII 56 (24): '8'
    rom[ 768] = 16'b0000000000000000;
    rom[ 769] = 16'b0000000000000000;
    rom[ 770] = 16'b0000000000000000;
    rom[ 771] = 16'b0000000000000000;
    rom[ 772] = 16'b0000000000000000;
    rom[ 773] = 16'b0000000000000000;
    rom[ 774] = 16'b0000000000000000;
    rom[ 775] = 16'b0000000000000000;
    rom[ 776] = 16'b0000000000000000;
    rom[ 777] = 16'b0000111111000000;
    rom[ 778] = 16'b0001111111100000;
    rom[ 779] = 16'b0011100001110000;
    rom[ 780] = 16'b0011000000110000;
    rom[ 781] = 16'b0011000000110000;
    rom[ 782] = 16'b0001110011100000;
    rom[ 783] = 16'b0000111111000000;
    rom[ 784] = 16'b0000111111000000;
    rom[ 785] = 16'b0001110011100000;
    rom[ 786] = 16'b0011100001110000;
    rom[ 787] = 16'b0011000000110000;
    rom[ 788] = 16'b0011000000110000;
    rom[ 789] = 16'b0011100001110000;
    rom[ 790] = 16'b0001111111100000;
    rom[ 791] = 16'b0000111111000000;
    rom[ 792] = 16'b0000000000000000;
    rom[ 793] = 16'b0000000000000000;
    rom[ 794] = 16'b0000000000000000;
    rom[ 795] = 16'b0000000000000000;
    rom[ 796] = 16'b0000000000000000;
    rom[ 797] = 16'b0000000000000000;
    rom[ 798] = 16'b0000000000000000;
    rom[ 799] = 16'b0000000000000000;

    // ASCII 57 (25): '9'
    rom[ 800] = 16'b0000000000000000;
    rom[ 801] = 16'b0000000000000000;
    rom[ 802] = 16'b0000000000000000;
    rom[ 803] = 16'b0000000000000000;
    rom[ 804] = 16'b0000000000000000;
    rom[ 805] = 16'b0000000000000000;
    rom[ 806] = 16'b0000000000000000;
    rom[ 807] = 16'b0000000000000000;
    rom[ 808] = 16'b0000000000000000;
    rom[ 809] = 16'b0000011110000000;
    rom[ 810] = 16'b0001111111100000;
    rom[ 811] = 16'b0001100001100000;
    rom[ 812] = 16'b0011000000110000;
    rom[ 813] = 16'b0011000000110000;
    rom[ 814] = 16'b0011000000110000;
    rom[ 815] = 16'b0011100001110000;
    rom[ 816] = 16'b0001111111110000;
    rom[ 817] = 16'b0000111110110000;
    rom[ 818] = 16'b0000000000110000;
    rom[ 819] = 16'b0000000001100000;
    rom[ 820] = 16'b0000000001100000;
    rom[ 821] = 16'b0000000111000000;
    rom[ 822] = 16'b0001111110000000;
    rom[ 823] = 16'b0001111100000000;
    rom[ 824] = 16'b0000000000000000;
    rom[ 825] = 16'b0000000000000000;
    rom[ 826] = 16'b0000000000000000;
    rom[ 827] = 16'b0000000000000000;
    rom[ 828] = 16'b0000000000000000;
    rom[ 829] = 16'b0000000000000000;
    rom[ 830] = 16'b0000000000000000;
    rom[ 831] = 16'b0000000000000000;

    // ASCII 58 (26): ':'
    rom[ 832] = 16'b0000000000000000;
    rom[ 833] = 16'b0000000000000000;
    rom[ 834] = 16'b0000000000000000;
    rom[ 835] = 16'b0000000000000000;
    rom[ 836] = 16'b0000000000000000;
    rom[ 837] = 16'b0000000000000000;
    rom[ 838] = 16'b0000000000000000;
    rom[ 839] = 16'b0000000000000000;
    rom[ 840] = 16'b0000000000000000;
    rom[ 841] = 16'b0000000000000000;
    rom[ 842] = 16'b0000000000000000;
    rom[ 843] = 16'b0000000000000000;
    rom[ 844] = 16'b0000000000000000;
    rom[ 845] = 16'b0000000000000000;
    rom[ 846] = 16'b0000000100000000;
    rom[ 847] = 16'b0000001110000000;
    rom[ 848] = 16'b0000001110000000;
    rom[ 849] = 16'b0000000100000000;
    rom[ 850] = 16'b0000000000000000;
    rom[ 851] = 16'b0000000000000000;
    rom[ 852] = 16'b0000000000000000;
    rom[ 853] = 16'b0000000000000000;
    rom[ 854] = 16'b0000000100000000;
    rom[ 855] = 16'b0000001110000000;
    rom[ 856] = 16'b0000001110000000;
    rom[ 857] = 16'b0000000100000000;
    rom[ 858] = 16'b0000000000000000;
    rom[ 859] = 16'b0000000000000000;
    rom[ 860] = 16'b0000000000000000;
    rom[ 861] = 16'b0000000000000000;
    rom[ 862] = 16'b0000000000000000;
    rom[ 863] = 16'b0000000000000000;

    // ASCII 59 (27): ';'
    rom[ 864] = 16'b0000000000000000;
    rom[ 865] = 16'b0000000000000000;
    rom[ 866] = 16'b0000000000000000;
    rom[ 867] = 16'b0000000000000000;
    rom[ 868] = 16'b0000000000000000;
    rom[ 869] = 16'b0000000000000000;
    rom[ 870] = 16'b0000000000000000;
    rom[ 871] = 16'b0000000000000000;
    rom[ 872] = 16'b0000000000000000;
    rom[ 873] = 16'b0000000000000000;
    rom[ 874] = 16'b0000000000000000;
    rom[ 875] = 16'b0000000000000000;
    rom[ 876] = 16'b0000000100000000;
    rom[ 877] = 16'b0000001110000000;
    rom[ 878] = 16'b0000001110000000;
    rom[ 879] = 16'b0000000100000000;
    rom[ 880] = 16'b0000000000000000;
    rom[ 881] = 16'b0000000000000000;
    rom[ 882] = 16'b0000000000000000;
    rom[ 883] = 16'b0000000000000000;
    rom[ 884] = 16'b0000001110000000;
    rom[ 885] = 16'b0000001111000000;
    rom[ 886] = 16'b0000001111000000;
    rom[ 887] = 16'b0000000111000000;
    rom[ 888] = 16'b0000000111000000;
    rom[ 889] = 16'b0000001110000000;
    rom[ 890] = 16'b0000111100000000;
    rom[ 891] = 16'b0000111000000000;
    rom[ 892] = 16'b0000000000000000;
    rom[ 893] = 16'b0000000000000000;
    rom[ 894] = 16'b0000000000000000;
    rom[ 895] = 16'b0000000000000000;

    // ASCII 60 (28): '<'
    rom[ 896] = 16'b0000000000000000;
    rom[ 897] = 16'b0000000000000000;
    rom[ 898] = 16'b0000000000000000;
    rom[ 899] = 16'b0000000000000000;
    rom[ 900] = 16'b0000000000000000;
    rom[ 901] = 16'b0000000000000000;
    rom[ 902] = 16'b0000000000000000;
    rom[ 903] = 16'b0000000000000000;
    rom[ 904] = 16'b0000000000000000;
    rom[ 905] = 16'b0000000000000000;
    rom[ 906] = 16'b0000000000000000;
    rom[ 907] = 16'b0000000000000000;
    rom[ 908] = 16'b0000000000100000;
    rom[ 909] = 16'b0000000001110000;
    rom[ 910] = 16'b0000000011100000;
    rom[ 911] = 16'b0000000110000000;
    rom[ 912] = 16'b0000011100000000;
    rom[ 913] = 16'b0000111000000000;
    rom[ 914] = 16'b0001110000000000;
    rom[ 915] = 16'b0000111000000000;
    rom[ 916] = 16'b0000011100000000;
    rom[ 917] = 16'b0000000110000000;
    rom[ 918] = 16'b0000000011100000;
    rom[ 919] = 16'b0000000001110000;
    rom[ 920] = 16'b0000000000100000;
    rom[ 921] = 16'b0000000000000000;
    rom[ 922] = 16'b0000000000000000;
    rom[ 923] = 16'b0000000000000000;
    rom[ 924] = 16'b0000000000000000;
    rom[ 925] = 16'b0000000000000000;
    rom[ 926] = 16'b0000000000000000;
    rom[ 927] = 16'b0000000000000000;

    // ASCII 61 (29): '='
    rom[ 928] = 16'b0000000000000000;
    rom[ 929] = 16'b0000000000000000;
    rom[ 930] = 16'b0000000000000000;
    rom[ 931] = 16'b0000000000000000;
    rom[ 932] = 16'b0000000000000000;
    rom[ 933] = 16'b0000000000000000;
    rom[ 934] = 16'b0000000000000000;
    rom[ 935] = 16'b0000000000000000;
    rom[ 936] = 16'b0000000000000000;
    rom[ 937] = 16'b0000000000000000;
    rom[ 938] = 16'b0000000000000000;
    rom[ 939] = 16'b0000000000000000;
    rom[ 940] = 16'b0000000000000000;
    rom[ 941] = 16'b0000000000000000;
    rom[ 942] = 16'b0000000000000000;
    rom[ 943] = 16'b0000000000000000;
    rom[ 944] = 16'b0000000000000000;
    rom[ 945] = 16'b0001111111111000;
    rom[ 946] = 16'b0001111111111000;
    rom[ 947] = 16'b0000000000000000;
    rom[ 948] = 16'b0000000000000000;
    rom[ 949] = 16'b0001111111111000;
    rom[ 950] = 16'b0001111111111000;
    rom[ 951] = 16'b0000000000000000;
    rom[ 952] = 16'b0000000000000000;
    rom[ 953] = 16'b0000000000000000;
    rom[ 954] = 16'b0000000000000000;
    rom[ 955] = 16'b0000000000000000;
    rom[ 956] = 16'b0000000000000000;
    rom[ 957] = 16'b0000000000000000;
    rom[ 958] = 16'b0000000000000000;
    rom[ 959] = 16'b0000000000000000;

    // ASCII 62 (30): '>'
    rom[ 960] = 16'b0000000000000000;
    rom[ 961] = 16'b0000000000000000;
    rom[ 962] = 16'b0000000000000000;
    rom[ 963] = 16'b0000000000000000;
    rom[ 964] = 16'b0000000000000000;
    rom[ 965] = 16'b0000000000000000;
    rom[ 966] = 16'b0000000000000000;
    rom[ 967] = 16'b0000000000000000;
    rom[ 968] = 16'b0000000000000000;
    rom[ 969] = 16'b0000000000000000;
    rom[ 970] = 16'b0000000000000000;
    rom[ 971] = 16'b0000000000000000;
    rom[ 972] = 16'b0000100000000000;
    rom[ 973] = 16'b0001110000000000;
    rom[ 974] = 16'b0000111000000000;
    rom[ 975] = 16'b0000001100000000;
    rom[ 976] = 16'b0000000111000000;
    rom[ 977] = 16'b0000000011100000;
    rom[ 978] = 16'b0000000001110000;
    rom[ 979] = 16'b0000000011100000;
    rom[ 980] = 16'b0000000111000000;
    rom[ 981] = 16'b0000001100000000;
    rom[ 982] = 16'b0000111000000000;
    rom[ 983] = 16'b0001110000000000;
    rom[ 984] = 16'b0000100000000000;
    rom[ 985] = 16'b0000000000000000;
    rom[ 986] = 16'b0000000000000000;
    rom[ 987] = 16'b0000000000000000;
    rom[ 988] = 16'b0000000000000000;
    rom[ 989] = 16'b0000000000000000;
    rom[ 990] = 16'b0000000000000000;
    rom[ 991] = 16'b0000000000000000;

    // ASCII 63 (31): '?'
    rom[ 992] = 16'b0000000000000000;
    rom[ 993] = 16'b0000000000000000;
    rom[ 994] = 16'b0000000000000000;
    rom[ 995] = 16'b0000000000000000;
    rom[ 996] = 16'b0000000000000000;
    rom[ 997] = 16'b0000000000000000;
    rom[ 998] = 16'b0000011100000000;
    rom[ 999] = 16'b0000011111000000;
    rom[1000] = 16'b0000000011100000;
    rom[1001] = 16'b0000000001110000;
    rom[1002] = 16'b0000000000110000;
    rom[1003] = 16'b0000000000110000;
    rom[1004] = 16'b0000000000110000;
    rom[1005] = 16'b0000000001110000;
    rom[1006] = 16'b0000000111100000;
    rom[1007] = 16'b0000000111000000;
    rom[1008] = 16'b0000000110000000;
    rom[1009] = 16'b0000000110000000;
    rom[1010] = 16'b0000000000000000;
    rom[1011] = 16'b0000000000000000;
    rom[1012] = 16'b0000001110000000;
    rom[1013] = 16'b0000001110000000;
    rom[1014] = 16'b0000001110000000;
    rom[1015] = 16'b0000000000000000;
    rom[1016] = 16'b0000000000000000;
    rom[1017] = 16'b0000000000000000;
    rom[1018] = 16'b0000000000000000;
    rom[1019] = 16'b0000000000000000;
    rom[1020] = 16'b0000000000000000;
    rom[1021] = 16'b0000000000000000;
    rom[1022] = 16'b0000000000000000;
    rom[1023] = 16'b0000000000000000;

    // ASCII 64 (32): '@'
    rom[1024] = 16'b0000000000000000;
    rom[1025] = 16'b0000000000000000;
    rom[1026] = 16'b0000000000000000;
    rom[1027] = 16'b0000000000000000;
    rom[1028] = 16'b0000011111000000;
    rom[1029] = 16'b0000110001100000;
    rom[1030] = 16'b0001100000110000;
    rom[1031] = 16'b0011000000110000;
    rom[1032] = 16'b0011000000011000;
    rom[1033] = 16'b0110000000011000;
    rom[1034] = 16'b0110001111011000;
    rom[1035] = 16'b0110011111011000;
    rom[1036] = 16'b1100011011011000;
    rom[1037] = 16'b1100110011011000;
    rom[1038] = 16'b1100110010011000;
    rom[1039] = 16'b1100110110011000;
    rom[1040] = 16'b1100110110011000;
    rom[1041] = 16'b1100110110011000;
    rom[1042] = 16'b1100110110110000;
    rom[1043] = 16'b1100111011110000;
    rom[1044] = 16'b1100011011100000;
    rom[1045] = 16'b0110000000000000;
    rom[1046] = 16'b0110000000000000;
    rom[1047] = 16'b0110000000000000;
    rom[1048] = 16'b0011100001000000;
    rom[1049] = 16'b0000111110000000;
    rom[1050] = 16'b0000000000000000;
    rom[1051] = 16'b0000000000000000;
    rom[1052] = 16'b0000000000000000;
    rom[1053] = 16'b0000000000000000;
    rom[1054] = 16'b0000000000000000;
    rom[1055] = 16'b0000000000000000;

    // ASCII 65 (33): 'A'
    rom[1056] = 16'b0000000000000000;
    rom[1057] = 16'b0000000000000000;
    rom[1058] = 16'b0000000000000000;
    rom[1059] = 16'b0000000000000000;
    rom[1060] = 16'b0000000000000000;
    rom[1061] = 16'b0000000000000000;
    rom[1062] = 16'b0000000000000000;
    rom[1063] = 16'b0000000000000000;
    rom[1064] = 16'b0000000000000000;
    rom[1065] = 16'b0000001110000000;
    rom[1066] = 16'b0000001011000000;
    rom[1067] = 16'b0000011011000000;
    rom[1068] = 16'b0000011011000000;
    rom[1069] = 16'b0000011001100000;
    rom[1070] = 16'b0000110001100000;
    rom[1071] = 16'b0000110001100000;
    rom[1072] = 16'b0000110000110000;
    rom[1073] = 16'b0000100000110000;
    rom[1074] = 16'b0001100000110000;
    rom[1075] = 16'b0001111111111000;
    rom[1076] = 16'b0001111111111000;
    rom[1077] = 16'b0011000000011100;
    rom[1078] = 16'b0011000000001100;
    rom[1079] = 16'b0011000000001100;
    rom[1080] = 16'b0000000000000000;
    rom[1081] = 16'b0000000000000000;
    rom[1082] = 16'b0000000000000000;
    rom[1083] = 16'b0000000000000000;
    rom[1084] = 16'b0000000000000000;
    rom[1085] = 16'b0000000000000000;
    rom[1086] = 16'b0000000000000000;
    rom[1087] = 16'b0000000000000000;

    // ASCII 66 (34): 'B'
    rom[1088] = 16'b0000000000000000;
    rom[1089] = 16'b0000000000000000;
    rom[1090] = 16'b0000000000000000;
    rom[1091] = 16'b0000000000000000;
    rom[1092] = 16'b0000000000000000;
    rom[1093] = 16'b0000000000000000;
    rom[1094] = 16'b0000000000000000;
    rom[1095] = 16'b0000000000000000;
    rom[1096] = 16'b0000000000000000;
    rom[1097] = 16'b0001111111000000;
    rom[1098] = 16'b0001111111100000;
    rom[1099] = 16'b0001100001110000;
    rom[1100] = 16'b0001100000110000;
    rom[1101] = 16'b0001100000110000;
    rom[1102] = 16'b0001100001100000;
    rom[1103] = 16'b0001111111000000;
    rom[1104] = 16'b0001111111110000;
    rom[1105] = 16'b0001100000110000;
    rom[1106] = 16'b0001100000011000;
    rom[1107] = 16'b0001100000011000;
    rom[1108] = 16'b0001100000011000;
    rom[1109] = 16'b0001100000110000;
    rom[1110] = 16'b0001111111110000;
    rom[1111] = 16'b0001111111000000;
    rom[1112] = 16'b0000000000000000;
    rom[1113] = 16'b0000000000000000;
    rom[1114] = 16'b0000000000000000;
    rom[1115] = 16'b0000000000000000;
    rom[1116] = 16'b0000000000000000;
    rom[1117] = 16'b0000000000000000;
    rom[1118] = 16'b0000000000000000;
    rom[1119] = 16'b0000000000000000;

    // ASCII 67 (35): 'C'
    rom[1120] = 16'b0000000000000000;
    rom[1121] = 16'b0000000000000000;
    rom[1122] = 16'b0000000000000000;
    rom[1123] = 16'b0000000000000000;
    rom[1124] = 16'b0000000000000000;
    rom[1125] = 16'b0000000000000000;
    rom[1126] = 16'b0000000000000000;
    rom[1127] = 16'b0000000000000000;
    rom[1128] = 16'b0000000000000000;
    rom[1129] = 16'b0000001111100000;
    rom[1130] = 16'b0000111111110000;
    rom[1131] = 16'b0001110000010000;
    rom[1132] = 16'b0001100000000000;
    rom[1133] = 16'b0011100000000000;
    rom[1134] = 16'b0011000000000000;
    rom[1135] = 16'b0011000000000000;
    rom[1136] = 16'b0011000000000000;
    rom[1137] = 16'b0011000000000000;
    rom[1138] = 16'b0011000000000000;
    rom[1139] = 16'b0011100000000000;
    rom[1140] = 16'b0001100000000000;
    rom[1141] = 16'b0001110000010000;
    rom[1142] = 16'b0000111111110000;
    rom[1143] = 16'b0000011111100000;
    rom[1144] = 16'b0000000000000000;
    rom[1145] = 16'b0000000000000000;
    rom[1146] = 16'b0000000000000000;
    rom[1147] = 16'b0000000000000000;
    rom[1148] = 16'b0000000000000000;
    rom[1149] = 16'b0000000000000000;
    rom[1150] = 16'b0000000000000000;
    rom[1151] = 16'b0000000000000000;

    // ASCII 68 (36): 'D'
    rom[1152] = 16'b0000000000000000;
    rom[1153] = 16'b0000000000000000;
    rom[1154] = 16'b0000000000000000;
    rom[1155] = 16'b0000000000000000;
    rom[1156] = 16'b0000000000000000;
    rom[1157] = 16'b0000000000000000;
    rom[1158] = 16'b0000000000000000;
    rom[1159] = 16'b0000000000000000;
    rom[1160] = 16'b0000000000000000;
    rom[1161] = 16'b0011111110000000;
    rom[1162] = 16'b0011111111100000;
    rom[1163] = 16'b0011000001110000;
    rom[1164] = 16'b0011000000110000;
    rom[1165] = 16'b0011000000011000;
    rom[1166] = 16'b0011000000011000;
    rom[1167] = 16'b0011000000011000;
    rom[1168] = 16'b0011000000011000;
    rom[1169] = 16'b0011000000011000;
    rom[1170] = 16'b0011000000011000;
    rom[1171] = 16'b0011000000111000;
    rom[1172] = 16'b0011000000110000;
    rom[1173] = 16'b0011000011110000;
    rom[1174] = 16'b0011111111100000;
    rom[1175] = 16'b0011111110000000;
    rom[1176] = 16'b0000000000000000;
    rom[1177] = 16'b0000000000000000;
    rom[1178] = 16'b0000000000000000;
    rom[1179] = 16'b0000000000000000;
    rom[1180] = 16'b0000000000000000;
    rom[1181] = 16'b0000000000000000;
    rom[1182] = 16'b0000000000000000;
    rom[1183] = 16'b0000000000000000;

    // ASCII 69 (37): 'E'
    rom[1184] = 16'b0000000000000000;
    rom[1185] = 16'b0000000000000000;
    rom[1186] = 16'b0000000000000000;
    rom[1187] = 16'b0000000000000000;
    rom[1188] = 16'b0000000000000000;
    rom[1189] = 16'b0000000000000000;
    rom[1190] = 16'b0000000000000000;
    rom[1191] = 16'b0000000000000000;
    rom[1192] = 16'b0000000000000000;
    rom[1193] = 16'b0001111111110000;
    rom[1194] = 16'b0001111111110000;
    rom[1195] = 16'b0001100000000000;
    rom[1196] = 16'b0001100000000000;
    rom[1197] = 16'b0001100000000000;
    rom[1198] = 16'b0001100000000000;
    rom[1199] = 16'b0001111111110000;
    rom[1200] = 16'b0001111111110000;
    rom[1201] = 16'b0001100000000000;
    rom[1202] = 16'b0001100000000000;
    rom[1203] = 16'b0001100000000000;
    rom[1204] = 16'b0001100000000000;
    rom[1205] = 16'b0001100000000000;
    rom[1206] = 16'b0001111111110000;
    rom[1207] = 16'b0001111111110000;
    rom[1208] = 16'b0000000000000000;
    rom[1209] = 16'b0000000000000000;
    rom[1210] = 16'b0000000000000000;
    rom[1211] = 16'b0000000000000000;
    rom[1212] = 16'b0000000000000000;
    rom[1213] = 16'b0000000000000000;
    rom[1214] = 16'b0000000000000000;
    rom[1215] = 16'b0000000000000000;

    // ASCII 70 (38): 'F'
    rom[1216] = 16'b0000000000000000;
    rom[1217] = 16'b0000000000000000;
    rom[1218] = 16'b0000000000000000;
    rom[1219] = 16'b0000000000000000;
    rom[1220] = 16'b0000000000000000;
    rom[1221] = 16'b0000000000000000;
    rom[1222] = 16'b0000000000000000;
    rom[1223] = 16'b0000000000000000;
    rom[1224] = 16'b0000000000000000;
    rom[1225] = 16'b0001111111110000;
    rom[1226] = 16'b0001111111110000;
    rom[1227] = 16'b0001100000000000;
    rom[1228] = 16'b0001100000000000;
    rom[1229] = 16'b0001100000000000;
    rom[1230] = 16'b0001100000000000;
    rom[1231] = 16'b0001111111110000;
    rom[1232] = 16'b0001111111110000;
    rom[1233] = 16'b0001100000000000;
    rom[1234] = 16'b0001100000000000;
    rom[1235] = 16'b0001100000000000;
    rom[1236] = 16'b0001100000000000;
    rom[1237] = 16'b0001100000000000;
    rom[1238] = 16'b0001100000000000;
    rom[1239] = 16'b0001100000000000;
    rom[1240] = 16'b0000000000000000;
    rom[1241] = 16'b0000000000000000;
    rom[1242] = 16'b0000000000000000;
    rom[1243] = 16'b0000000000000000;
    rom[1244] = 16'b0000000000000000;
    rom[1245] = 16'b0000000000000000;
    rom[1246] = 16'b0000000000000000;
    rom[1247] = 16'b0000000000000000;

    // ASCII 71 (39): 'G'
    rom[1248] = 16'b0000000000000000;
    rom[1249] = 16'b0000000000000000;
    rom[1250] = 16'b0000000000000000;
    rom[1251] = 16'b0000000000000000;
    rom[1252] = 16'b0000000000000000;
    rom[1253] = 16'b0000000000000000;
    rom[1254] = 16'b0000000000000000;
    rom[1255] = 16'b0000000000000000;
    rom[1256] = 16'b0000000000000000;
    rom[1257] = 16'b0000001111110000;
    rom[1258] = 16'b0000011111111000;
    rom[1259] = 16'b0000111000001000;
    rom[1260] = 16'b0001100000000000;
    rom[1261] = 16'b0011100000000000;
    rom[1262] = 16'b0011000000000000;
    rom[1263] = 16'b0011000011111000;
    rom[1264] = 16'b0011000011111000;
    rom[1265] = 16'b0011000000011000;
    rom[1266] = 16'b0011000000011000;
    rom[1267] = 16'b0011100000011000;
    rom[1268] = 16'b0001100000011000;
    rom[1269] = 16'b0001110000011000;
    rom[1270] = 16'b0000111111111000;
    rom[1271] = 16'b0000001111110000;
    rom[1272] = 16'b0000000000000000;
    rom[1273] = 16'b0000000000000000;
    rom[1274] = 16'b0000000000000000;
    rom[1275] = 16'b0000000000000000;
    rom[1276] = 16'b0000000000000000;
    rom[1277] = 16'b0000000000000000;
    rom[1278] = 16'b0000000000000000;
    rom[1279] = 16'b0000000000000000;

    // ASCII 72 (40): 'H'
    rom[1280] = 16'b0000000000000000;
    rom[1281] = 16'b0000000000000000;
    rom[1282] = 16'b0000000000000000;
    rom[1283] = 16'b0000000000000000;
    rom[1284] = 16'b0000000000000000;
    rom[1285] = 16'b0000000000000000;
    rom[1286] = 16'b0000000000000000;
    rom[1287] = 16'b0000000000000000;
    rom[1288] = 16'b0000000000000000;
    rom[1289] = 16'b0011000000011000;
    rom[1290] = 16'b0011000000011000;
    rom[1291] = 16'b0011000000011000;
    rom[1292] = 16'b0011000000011000;
    rom[1293] = 16'b0011000000011000;
    rom[1294] = 16'b0011000000011000;
    rom[1295] = 16'b0011111111111000;
    rom[1296] = 16'b0011111111111000;
    rom[1297] = 16'b0011000000011000;
    rom[1298] = 16'b0011000000011000;
    rom[1299] = 16'b0011000000011000;
    rom[1300] = 16'b0011000000011000;
    rom[1301] = 16'b0011000000011000;
    rom[1302] = 16'b0011000000011000;
    rom[1303] = 16'b0011000000011000;
    rom[1304] = 16'b0000000000000000;
    rom[1305] = 16'b0000000000000000;
    rom[1306] = 16'b0000000000000000;
    rom[1307] = 16'b0000000000000000;
    rom[1308] = 16'b0000000000000000;
    rom[1309] = 16'b0000000000000000;
    rom[1310] = 16'b0000000000000000;
    rom[1311] = 16'b0000000000000000;

    // ASCII 73 (41): 'I'
    rom[1312] = 16'b0000000000000000;
    rom[1313] = 16'b0000000000000000;
    rom[1314] = 16'b0000000000000000;
    rom[1315] = 16'b0000000000000000;
    rom[1316] = 16'b0000000000000000;
    rom[1317] = 16'b0000000000000000;
    rom[1318] = 16'b0000000000000000;
    rom[1319] = 16'b0000000000000000;
    rom[1320] = 16'b0000000000000000;
    rom[1321] = 16'b0001111111111000;
    rom[1322] = 16'b0001111111111000;
    rom[1323] = 16'b0000000110000000;
    rom[1324] = 16'b0000000110000000;
    rom[1325] = 16'b0000000110000000;
    rom[1326] = 16'b0000000110000000;
    rom[1327] = 16'b0000000110000000;
    rom[1328] = 16'b0000000110000000;
    rom[1329] = 16'b0000000110000000;
    rom[1330] = 16'b0000000110000000;
    rom[1331] = 16'b0000000110000000;
    rom[1332] = 16'b0000000110000000;
    rom[1333] = 16'b0000000110000000;
    rom[1334] = 16'b0001111111111000;
    rom[1335] = 16'b0001111111111000;
    rom[1336] = 16'b0000000000000000;
    rom[1337] = 16'b0000000000000000;
    rom[1338] = 16'b0000000000000000;
    rom[1339] = 16'b0000000000000000;
    rom[1340] = 16'b0000000000000000;
    rom[1341] = 16'b0000000000000000;
    rom[1342] = 16'b0000000000000000;
    rom[1343] = 16'b0000000000000000;

    // ASCII 74 (42): 'J'
    rom[1344] = 16'b0000000000000000;
    rom[1345] = 16'b0000000000000000;
    rom[1346] = 16'b0000000000000000;
    rom[1347] = 16'b0000000000000000;
    rom[1348] = 16'b0000000000000000;
    rom[1349] = 16'b0000000000000000;
    rom[1350] = 16'b0000000000000000;
    rom[1351] = 16'b0000000000000000;
    rom[1352] = 16'b0000000000000000;
    rom[1353] = 16'b0001111111100000;
    rom[1354] = 16'b0001111111100000;
    rom[1355] = 16'b0000000001100000;
    rom[1356] = 16'b0000000001100000;
    rom[1357] = 16'b0000000001100000;
    rom[1358] = 16'b0000000001100000;
    rom[1359] = 16'b0000000001100000;
    rom[1360] = 16'b0000000001100000;
    rom[1361] = 16'b0000000001100000;
    rom[1362] = 16'b0000000001100000;
    rom[1363] = 16'b0000000001100000;
    rom[1364] = 16'b0000000001100000;
    rom[1365] = 16'b0001000011100000;
    rom[1366] = 16'b0001111111000000;
    rom[1367] = 16'b0000111110000000;
    rom[1368] = 16'b0000000000000000;
    rom[1369] = 16'b0000000000000000;
    rom[1370] = 16'b0000000000000000;
    rom[1371] = 16'b0000000000000000;
    rom[1372] = 16'b0000000000000000;
    rom[1373] = 16'b0000000000000000;
    rom[1374] = 16'b0000000000000000;
    rom[1375] = 16'b0000000000000000;

    // ASCII 75 (43): 'K'
    rom[1376] = 16'b0000000000000000;
    rom[1377] = 16'b0000000000000000;
    rom[1378] = 16'b0000000000000000;
    rom[1379] = 16'b0000000000000000;
    rom[1380] = 16'b0000000000000000;
    rom[1381] = 16'b0000000000000000;
    rom[1382] = 16'b0000000000000000;
    rom[1383] = 16'b0000000000000000;
    rom[1384] = 16'b0000000000000000;
    rom[1385] = 16'b0001100000011000;
    rom[1386] = 16'b0001100000110000;
    rom[1387] = 16'b0001100001100000;
    rom[1388] = 16'b0001100011000000;
    rom[1389] = 16'b0001100111000000;
    rom[1390] = 16'b0001100110000000;
    rom[1391] = 16'b0001101100000000;
    rom[1392] = 16'b0001111000000000;
    rom[1393] = 16'b0001101100000000;
    rom[1394] = 16'b0001100110000000;
    rom[1395] = 16'b0001100111000000;
    rom[1396] = 16'b0001100011100000;
    rom[1397] = 16'b0001100001100000;
    rom[1398] = 16'b0001100000110000;
    rom[1399] = 16'b0001100000011000;
    rom[1400] = 16'b0000000000000000;
    rom[1401] = 16'b0000000000000000;
    rom[1402] = 16'b0000000000000000;
    rom[1403] = 16'b0000000000000000;
    rom[1404] = 16'b0000000000000000;
    rom[1405] = 16'b0000000000000000;
    rom[1406] = 16'b0000000000000000;
    rom[1407] = 16'b0000000000000000;

    // ASCII 76 (44): 'L'
    rom[1408] = 16'b0000000000000000;
    rom[1409] = 16'b0000000000000000;
    rom[1410] = 16'b0000000000000000;
    rom[1411] = 16'b0000000000000000;
    rom[1412] = 16'b0000000000000000;
    rom[1413] = 16'b0000000000000000;
    rom[1414] = 16'b0000000000000000;
    rom[1415] = 16'b0000000000000000;
    rom[1416] = 16'b0000000000000000;
    rom[1417] = 16'b0000110000000000;
    rom[1418] = 16'b0000110000000000;
    rom[1419] = 16'b0000110000000000;
    rom[1420] = 16'b0000110000000000;
    rom[1421] = 16'b0000110000000000;
    rom[1422] = 16'b0000110000000000;
    rom[1423] = 16'b0000110000000000;
    rom[1424] = 16'b0000110000000000;
    rom[1425] = 16'b0000110000000000;
    rom[1426] = 16'b0000110000000000;
    rom[1427] = 16'b0000110000000000;
    rom[1428] = 16'b0000110000000000;
    rom[1429] = 16'b0000110000000000;
    rom[1430] = 16'b0000111111111000;
    rom[1431] = 16'b0000111111111000;
    rom[1432] = 16'b0000000000000000;
    rom[1433] = 16'b0000000000000000;
    rom[1434] = 16'b0000000000000000;
    rom[1435] = 16'b0000000000000000;
    rom[1436] = 16'b0000000000000000;
    rom[1437] = 16'b0000000000000000;
    rom[1438] = 16'b0000000000000000;
    rom[1439] = 16'b0000000000000000;

    // ASCII 77 (45): 'M'
    rom[1440] = 16'b0000000000000000;
    rom[1441] = 16'b0000000000000000;
    rom[1442] = 16'b0000000000000000;
    rom[1443] = 16'b0000000000000000;
    rom[1444] = 16'b0000000000000000;
    rom[1445] = 16'b0000000000000000;
    rom[1446] = 16'b0000000000000000;
    rom[1447] = 16'b0000000000000000;
    rom[1448] = 16'b0000000000000000;
    rom[1449] = 16'b0011100000111000;
    rom[1450] = 16'b0011100000111000;
    rom[1451] = 16'b0011100000111000;
    rom[1452] = 16'b0011110001111000;
    rom[1453] = 16'b0011010001011000;
    rom[1454] = 16'b0011011011011000;
    rom[1455] = 16'b0011011011011000;
    rom[1456] = 16'b0011001010011000;
    rom[1457] = 16'b0011001110011000;
    rom[1458] = 16'b0011001100011000;
    rom[1459] = 16'b0011000000011000;
    rom[1460] = 16'b0011000000011000;
    rom[1461] = 16'b0011000000011000;
    rom[1462] = 16'b0011000000011100;
    rom[1463] = 16'b0011000000011100;
    rom[1464] = 16'b0000000000000000;
    rom[1465] = 16'b0000000000000000;
    rom[1466] = 16'b0000000000000000;
    rom[1467] = 16'b0000000000000000;
    rom[1468] = 16'b0000000000000000;
    rom[1469] = 16'b0000000000000000;
    rom[1470] = 16'b0000000000000000;
    rom[1471] = 16'b0000000000000000;

    // ASCII 78 (46): 'N'
    rom[1472] = 16'b0000000000000000;
    rom[1473] = 16'b0000000000000000;
    rom[1474] = 16'b0000000000000000;
    rom[1475] = 16'b0000000000000000;
    rom[1476] = 16'b0000000000000000;
    rom[1477] = 16'b0000000000000000;
    rom[1478] = 16'b0000000000000000;
    rom[1479] = 16'b0000000000000000;
    rom[1480] = 16'b0000000000000000;
    rom[1481] = 16'b0011100000011000;
    rom[1482] = 16'b0011110000011000;
    rom[1483] = 16'b0011110000011000;
    rom[1484] = 16'b0011011000011000;
    rom[1485] = 16'b0011011000011000;
    rom[1486] = 16'b0011001000011000;
    rom[1487] = 16'b0011001100011000;
    rom[1488] = 16'b0011000100011000;
    rom[1489] = 16'b0011000110011000;
    rom[1490] = 16'b0011000110011000;
    rom[1491] = 16'b0011000011011000;
    rom[1492] = 16'b0011000011011000;
    rom[1493] = 16'b0011000001111000;
    rom[1494] = 16'b0011000001111000;
    rom[1495] = 16'b0011000000111000;
    rom[1496] = 16'b0000000000000000;
    rom[1497] = 16'b0000000000000000;
    rom[1498] = 16'b0000000000000000;
    rom[1499] = 16'b0000000000000000;
    rom[1500] = 16'b0000000000000000;
    rom[1501] = 16'b0000000000000000;
    rom[1502] = 16'b0000000000000000;
    rom[1503] = 16'b0000000000000000;

    // ASCII 79 (47): 'O'
    rom[1504] = 16'b0000000000000000;
    rom[1505] = 16'b0000000000000000;
    rom[1506] = 16'b0000000000000000;
    rom[1507] = 16'b0000000000000000;
    rom[1508] = 16'b0000000000000000;
    rom[1509] = 16'b0000000000000000;
    rom[1510] = 16'b0000000000000000;
    rom[1511] = 16'b0000000000000000;
    rom[1512] = 16'b0000000000000000;
    rom[1513] = 16'b0000001111100000;
    rom[1514] = 16'b0000111111110000;
    rom[1515] = 16'b0001110000111000;
    rom[1516] = 16'b0001100000011000;
    rom[1517] = 16'b0011000000001100;
    rom[1518] = 16'b0011000000001100;
    rom[1519] = 16'b0011000000001100;
    rom[1520] = 16'b0011000000001100;
    rom[1521] = 16'b0011000000001100;
    rom[1522] = 16'b0011000000001100;
    rom[1523] = 16'b0011000000011100;
    rom[1524] = 16'b0001100000011000;
    rom[1525] = 16'b0001110000111000;
    rom[1526] = 16'b0000111111110000;
    rom[1527] = 16'b0000011111000000;
    rom[1528] = 16'b0000000000000000;
    rom[1529] = 16'b0000000000000000;
    rom[1530] = 16'b0000000000000000;
    rom[1531] = 16'b0000000000000000;
    rom[1532] = 16'b0000000000000000;
    rom[1533] = 16'b0000000000000000;
    rom[1534] = 16'b0000000000000000;
    rom[1535] = 16'b0000000000000000;

    // ASCII 80 (48): 'P'
    rom[1536] = 16'b0000000000000000;
    rom[1537] = 16'b0000000000000000;
    rom[1538] = 16'b0000000000000000;
    rom[1539] = 16'b0000000000000000;
    rom[1540] = 16'b0000000000000000;
    rom[1541] = 16'b0000000000000000;
    rom[1542] = 16'b0000000000000000;
    rom[1543] = 16'b0000000000000000;
    rom[1544] = 16'b0000000000000000;
    rom[1545] = 16'b0001111111000000;
    rom[1546] = 16'b0001111111110000;
    rom[1547] = 16'b0001100000111000;
    rom[1548] = 16'b0001100000011000;
    rom[1549] = 16'b0001100000011000;
    rom[1550] = 16'b0001100000011000;
    rom[1551] = 16'b0001100000011000;
    rom[1552] = 16'b0001100001110000;
    rom[1553] = 16'b0001111111100000;
    rom[1554] = 16'b0001111111000000;
    rom[1555] = 16'b0001100000000000;
    rom[1556] = 16'b0001100000000000;
    rom[1557] = 16'b0001100000000000;
    rom[1558] = 16'b0001100000000000;
    rom[1559] = 16'b0001100000000000;
    rom[1560] = 16'b0000000000000000;
    rom[1561] = 16'b0000000000000000;
    rom[1562] = 16'b0000000000000000;
    rom[1563] = 16'b0000000000000000;
    rom[1564] = 16'b0000000000000000;
    rom[1565] = 16'b0000000000000000;
    rom[1566] = 16'b0000000000000000;
    rom[1567] = 16'b0000000000000000;

    // ASCII 81 (49): 'Q'
    rom[1568] = 16'b0000000000000000;
    rom[1569] = 16'b0000000000000000;
    rom[1570] = 16'b0000000000000000;
    rom[1571] = 16'b0000000000000000;
    rom[1572] = 16'b0000000000000000;
    rom[1573] = 16'b0000000000000000;
    rom[1574] = 16'b0000000000000000;
    rom[1575] = 16'b0000001111100000;
    rom[1576] = 16'b0000111111110000;
    rom[1577] = 16'b0001110000111000;
    rom[1578] = 16'b0001100000011000;
    rom[1579] = 16'b0011000000001100;
    rom[1580] = 16'b0011000000001100;
    rom[1581] = 16'b0011000000001100;
    rom[1582] = 16'b0011000000001100;
    rom[1583] = 16'b0011000000001100;
    rom[1584] = 16'b0011000000001100;
    rom[1585] = 16'b0011000000011100;
    rom[1586] = 16'b0001100000011000;
    rom[1587] = 16'b0001110000111000;
    rom[1588] = 16'b0000111111110000;
    rom[1589] = 16'b0000011111100000;
    rom[1590] = 16'b0000000110000000;
    rom[1591] = 16'b0000000111000110;
    rom[1592] = 16'b0000000011111110;
    rom[1593] = 16'b0000000001111000;
    rom[1594] = 16'b0000000000000000;
    rom[1595] = 16'b0000000000000000;
    rom[1596] = 16'b0000000000000000;
    rom[1597] = 16'b0000000000000000;
    rom[1598] = 16'b0000000000000000;
    rom[1599] = 16'b0000000000000000;

    // ASCII 82 (50): 'R'
    rom[1600] = 16'b0000000000000000;
    rom[1601] = 16'b0000000000000000;
    rom[1602] = 16'b0000000000000000;
    rom[1603] = 16'b0000000000000000;
    rom[1604] = 16'b0000000000000000;
    rom[1605] = 16'b0000000000000000;
    rom[1606] = 16'b0000000000000000;
    rom[1607] = 16'b0000000000000000;
    rom[1608] = 16'b0000000000000000;
    rom[1609] = 16'b0001111111000000;
    rom[1610] = 16'b0001111111100000;
    rom[1611] = 16'b0001100001110000;
    rom[1612] = 16'b0001100000110000;
    rom[1613] = 16'b0001100000110000;
    rom[1614] = 16'b0001100000110000;
    rom[1615] = 16'b0001100001100000;
    rom[1616] = 16'b0001111111100000;
    rom[1617] = 16'b0001111110000000;
    rom[1618] = 16'b0001100011000000;
    rom[1619] = 16'b0001100011100000;
    rom[1620] = 16'b0001100001100000;
    rom[1621] = 16'b0001100001110000;
    rom[1622] = 16'b0001100000110000;
    rom[1623] = 16'b0001100000111000;
    rom[1624] = 16'b0000000000000000;
    rom[1625] = 16'b0000000000000000;
    rom[1626] = 16'b0000000000000000;
    rom[1627] = 16'b0000000000000000;
    rom[1628] = 16'b0000000000000000;
    rom[1629] = 16'b0000000000000000;
    rom[1630] = 16'b0000000000000000;
    rom[1631] = 16'b0000000000000000;

    // ASCII 83 (51): 'S'
    rom[1632] = 16'b0000000000000000;
    rom[1633] = 16'b0000000000000000;
    rom[1634] = 16'b0000000000000000;
    rom[1635] = 16'b0000000000000000;
    rom[1636] = 16'b0000000000000000;
    rom[1637] = 16'b0000000000000000;
    rom[1638] = 16'b0000000000000000;
    rom[1639] = 16'b0000000000000000;
    rom[1640] = 16'b0000000000000000;
    rom[1641] = 16'b0000011111000000;
    rom[1642] = 16'b0001111111100000;
    rom[1643] = 16'b0011100000100000;
    rom[1644] = 16'b0011000000000000;
    rom[1645] = 16'b0011000000000000;
    rom[1646] = 16'b0011100000000000;
    rom[1647] = 16'b0001111000000000;
    rom[1648] = 16'b0000011111000000;
    rom[1649] = 16'b0000000111100000;
    rom[1650] = 16'b0000000001110000;
    rom[1651] = 16'b0000000000110000;
    rom[1652] = 16'b0000000000110000;
    rom[1653] = 16'b0010000001110000;
    rom[1654] = 16'b0011111111100000;
    rom[1655] = 16'b0001111110000000;
    rom[1656] = 16'b0000000000000000;
    rom[1657] = 16'b0000000000000000;
    rom[1658] = 16'b0000000000000000;
    rom[1659] = 16'b0000000000000000;
    rom[1660] = 16'b0000000000000000;
    rom[1661] = 16'b0000000000000000;
    rom[1662] = 16'b0000000000000000;
    rom[1663] = 16'b0000000000000000;

    // ASCII 84 (52): 'T'
    rom[1664] = 16'b0000000000000000;
    rom[1665] = 16'b0000000000000000;
    rom[1666] = 16'b0000000000000000;
    rom[1667] = 16'b0000000000000000;
    rom[1668] = 16'b0000000000000000;
    rom[1669] = 16'b0000000000000000;
    rom[1670] = 16'b0000000000000000;
    rom[1671] = 16'b0000000000000000;
    rom[1672] = 16'b0000000000000000;
    rom[1673] = 16'b0011111111111100;
    rom[1674] = 16'b0011111111111100;
    rom[1675] = 16'b0000000110000000;
    rom[1676] = 16'b0000000110000000;
    rom[1677] = 16'b0000000110000000;
    rom[1678] = 16'b0000000110000000;
    rom[1679] = 16'b0000000110000000;
    rom[1680] = 16'b0000000110000000;
    rom[1681] = 16'b0000000110000000;
    rom[1682] = 16'b0000000110000000;
    rom[1683] = 16'b0000000110000000;
    rom[1684] = 16'b0000000110000000;
    rom[1685] = 16'b0000000110000000;
    rom[1686] = 16'b0000000110000000;
    rom[1687] = 16'b0000000110000000;
    rom[1688] = 16'b0000000000000000;
    rom[1689] = 16'b0000000000000000;
    rom[1690] = 16'b0000000000000000;
    rom[1691] = 16'b0000000000000000;
    rom[1692] = 16'b0000000000000000;
    rom[1693] = 16'b0000000000000000;
    rom[1694] = 16'b0000000000000000;
    rom[1695] = 16'b0000000000000000;

    // ASCII 85 (53): 'U'
    rom[1696] = 16'b0000000000000000;
    rom[1697] = 16'b0000000000000000;
    rom[1698] = 16'b0000000000000000;
    rom[1699] = 16'b0000000000000000;
    rom[1700] = 16'b0000000000000000;
    rom[1701] = 16'b0000000000000000;
    rom[1702] = 16'b0000000000000000;
    rom[1703] = 16'b0000000000000000;
    rom[1704] = 16'b0000000000000000;
    rom[1705] = 16'b0011000000011000;
    rom[1706] = 16'b0011000000011000;
    rom[1707] = 16'b0011000000011000;
    rom[1708] = 16'b0011000000011000;
    rom[1709] = 16'b0011000000011000;
    rom[1710] = 16'b0011000000011000;
    rom[1711] = 16'b0011000000011000;
    rom[1712] = 16'b0011000000011000;
    rom[1713] = 16'b0011000000011000;
    rom[1714] = 16'b0011000000011000;
    rom[1715] = 16'b0011000000011000;
    rom[1716] = 16'b0011000000011000;
    rom[1717] = 16'b0011100000110000;
    rom[1718] = 16'b0001111111110000;
    rom[1719] = 16'b0000011111000000;
    rom[1720] = 16'b0000000000000000;
    rom[1721] = 16'b0000000000000000;
    rom[1722] = 16'b0000000000000000;
    rom[1723] = 16'b0000000000000000;
    rom[1724] = 16'b0000000000000000;
    rom[1725] = 16'b0000000000000000;
    rom[1726] = 16'b0000000000000000;
    rom[1727] = 16'b0000000000000000;

    // ASCII 86 (54): 'V'
    rom[1728] = 16'b0000000000000000;
    rom[1729] = 16'b0000000000000000;
    rom[1730] = 16'b0000000000000000;
    rom[1731] = 16'b0000000000000000;
    rom[1732] = 16'b0000000000000000;
    rom[1733] = 16'b0000000000000000;
    rom[1734] = 16'b0000000000000000;
    rom[1735] = 16'b0000000000000000;
    rom[1736] = 16'b0000000000000000;
    rom[1737] = 16'b1100000000011000;
    rom[1738] = 16'b1100000000011000;
    rom[1739] = 16'b1110000000111000;
    rom[1740] = 16'b0110000000110000;
    rom[1741] = 16'b0110000000110000;
    rom[1742] = 16'b0011000001100000;
    rom[1743] = 16'b0011000001100000;
    rom[1744] = 16'b0011100001100000;
    rom[1745] = 16'b0001100011000000;
    rom[1746] = 16'b0001100011000000;
    rom[1747] = 16'b0001110111000000;
    rom[1748] = 16'b0000110110000000;
    rom[1749] = 16'b0000110110000000;
    rom[1750] = 16'b0000111100000000;
    rom[1751] = 16'b0000011100000000;
    rom[1752] = 16'b0000000000000000;
    rom[1753] = 16'b0000000000000000;
    rom[1754] = 16'b0000000000000000;
    rom[1755] = 16'b0000000000000000;
    rom[1756] = 16'b0000000000000000;
    rom[1757] = 16'b0000000000000000;
    rom[1758] = 16'b0000000000000000;
    rom[1759] = 16'b0000000000000000;

    // ASCII 87 (55): 'W'
    rom[1760] = 16'b0000000000000000;
    rom[1761] = 16'b0000000000000000;
    rom[1762] = 16'b0000000000000000;
    rom[1763] = 16'b0000000000000000;
    rom[1764] = 16'b0000000000000000;
    rom[1765] = 16'b0000000000000000;
    rom[1766] = 16'b0000000000000000;
    rom[1767] = 16'b0000000000000000;
    rom[1768] = 16'b0000000000000000;
    rom[1769] = 16'b0011000000011000;
    rom[1770] = 16'b0011000000011000;
    rom[1771] = 16'b0011000000011000;
    rom[1772] = 16'b0011000000011000;
    rom[1773] = 16'b0011000000011000;
    rom[1774] = 16'b0011000100011000;
    rom[1775] = 16'b0011000110011000;
    rom[1776] = 16'b0011001010011000;
    rom[1777] = 16'b0011001010011000;
    rom[1778] = 16'b0011001010011000;
    rom[1779] = 16'b0001101011010000;
    rom[1780] = 16'b0001111011110000;
    rom[1781] = 16'b0001111011110000;
    rom[1782] = 16'b0001110001110000;
    rom[1783] = 16'b0001110001110000;
    rom[1784] = 16'b0000000000000000;
    rom[1785] = 16'b0000000000000000;
    rom[1786] = 16'b0000000000000000;
    rom[1787] = 16'b0000000000000000;
    rom[1788] = 16'b0000000000000000;
    rom[1789] = 16'b0000000000000000;
    rom[1790] = 16'b0000000000000000;
    rom[1791] = 16'b0000000000000000;

    // ASCII 88 (56): 'X'
    rom[1792] = 16'b0000000000000000;
    rom[1793] = 16'b0000000000000000;
    rom[1794] = 16'b0000000000000000;
    rom[1795] = 16'b0000000000000000;
    rom[1796] = 16'b0000000000000000;
    rom[1797] = 16'b0000000000000000;
    rom[1798] = 16'b0000000000000000;
    rom[1799] = 16'b0000000000000000;
    rom[1800] = 16'b0000000000000000;
    rom[1801] = 16'b0011100000011100;
    rom[1802] = 16'b0001100000011000;
    rom[1803] = 16'b0000110000110000;
    rom[1804] = 16'b0000111001110000;
    rom[1805] = 16'b0000011011100000;
    rom[1806] = 16'b0000011111000000;
    rom[1807] = 16'b0000001111000000;
    rom[1808] = 16'b0000001110000000;
    rom[1809] = 16'b0000001111000000;
    rom[1810] = 16'b0000011011100000;
    rom[1811] = 16'b0000111001100000;
    rom[1812] = 16'b0001110001110000;
    rom[1813] = 16'b0001100000110000;
    rom[1814] = 16'b0011100000111000;
    rom[1815] = 16'b0111000000011100;
    rom[1816] = 16'b0000000000000000;
    rom[1817] = 16'b0000000000000000;
    rom[1818] = 16'b0000000000000000;
    rom[1819] = 16'b0000000000000000;
    rom[1820] = 16'b0000000000000000;
    rom[1821] = 16'b0000000000000000;
    rom[1822] = 16'b0000000000000000;
    rom[1823] = 16'b0000000000000000;

    // ASCII 89 (57): 'Y'
    rom[1824] = 16'b0000000000000000;
    rom[1825] = 16'b0000000000000000;
    rom[1826] = 16'b0000000000000000;
    rom[1827] = 16'b0000000000000000;
    rom[1828] = 16'b0000000000000000;
    rom[1829] = 16'b0000000000000000;
    rom[1830] = 16'b0000000000000000;
    rom[1831] = 16'b0000000000000000;
    rom[1832] = 16'b0000000000000000;
    rom[1833] = 16'b1100000000001100;
    rom[1834] = 16'b0110000000011000;
    rom[1835] = 16'b0111000000111000;
    rom[1836] = 16'b0011000000110000;
    rom[1837] = 16'b0001100001100000;
    rom[1838] = 16'b0001110001100000;
    rom[1839] = 16'b0000110011000000;
    rom[1840] = 16'b0000111111000000;
    rom[1841] = 16'b0000011110000000;
    rom[1842] = 16'b0000001100000000;
    rom[1843] = 16'b0000001100000000;
    rom[1844] = 16'b0000001100000000;
    rom[1845] = 16'b0000001100000000;
    rom[1846] = 16'b0000001100000000;
    rom[1847] = 16'b0000001100000000;
    rom[1848] = 16'b0000000000000000;
    rom[1849] = 16'b0000000000000000;
    rom[1850] = 16'b0000000000000000;
    rom[1851] = 16'b0000000000000000;
    rom[1852] = 16'b0000000000000000;
    rom[1853] = 16'b0000000000000000;
    rom[1854] = 16'b0000000000000000;
    rom[1855] = 16'b0000000000000000;

    // ASCII 90 (58): 'Z'
    rom[1856] = 16'b0000000000000000;
    rom[1857] = 16'b0000000000000000;
    rom[1858] = 16'b0000000000000000;
    rom[1859] = 16'b0000000000000000;
    rom[1860] = 16'b0000000000000000;
    rom[1861] = 16'b0000000000000000;
    rom[1862] = 16'b0000000000000000;
    rom[1863] = 16'b0000000000000000;
    rom[1864] = 16'b0000000000000000;
    rom[1865] = 16'b0011111111110000;
    rom[1866] = 16'b0011111111110000;
    rom[1867] = 16'b0000000001100000;
    rom[1868] = 16'b0000000011100000;
    rom[1869] = 16'b0000000011000000;
    rom[1870] = 16'b0000000110000000;
    rom[1871] = 16'b0000000110000000;
    rom[1872] = 16'b0000001100000000;
    rom[1873] = 16'b0000011000000000;
    rom[1874] = 16'b0000011000000000;
    rom[1875] = 16'b0000110000000000;
    rom[1876] = 16'b0001110000000000;
    rom[1877] = 16'b0001100000000000;
    rom[1878] = 16'b0011111111111000;
    rom[1879] = 16'b0011111111111000;
    rom[1880] = 16'b0000000000000000;
    rom[1881] = 16'b0000000000000000;
    rom[1882] = 16'b0000000000000000;
    rom[1883] = 16'b0000000000000000;
    rom[1884] = 16'b0000000000000000;
    rom[1885] = 16'b0000000000000000;
    rom[1886] = 16'b0000000000000000;
    rom[1887] = 16'b0000000000000000;

    // ASCII 91 (59): '['
    rom[1888] = 16'b0000000000000000;
    rom[1889] = 16'b0000000000000000;
    rom[1890] = 16'b0000000000000000;
    rom[1891] = 16'b0000000000000000;
    rom[1892] = 16'b0000011111100000;
    rom[1893] = 16'b0000011111100000;
    rom[1894] = 16'b0000011000000000;
    rom[1895] = 16'b0000011000000000;
    rom[1896] = 16'b0000011000000000;
    rom[1897] = 16'b0000011000000000;
    rom[1898] = 16'b0000011000000000;
    rom[1899] = 16'b0000011000000000;
    rom[1900] = 16'b0000011000000000;
    rom[1901] = 16'b0000011000000000;
    rom[1902] = 16'b0000011000000000;
    rom[1903] = 16'b0000011000000000;
    rom[1904] = 16'b0000011000000000;
    rom[1905] = 16'b0000011000000000;
    rom[1906] = 16'b0000011000000000;
    rom[1907] = 16'b0000011000000000;
    rom[1908] = 16'b0000011000000000;
    rom[1909] = 16'b0000011000000000;
    rom[1910] = 16'b0000011000000000;
    rom[1911] = 16'b0000011000000000;
    rom[1912] = 16'b0000011111100000;
    rom[1913] = 16'b0000011111100000;
    rom[1914] = 16'b0000000000000000;
    rom[1915] = 16'b0000000000000000;
    rom[1916] = 16'b0000000000000000;
    rom[1917] = 16'b0000000000000000;
    rom[1918] = 16'b0000000000000000;
    rom[1919] = 16'b0000000000000000;

    // ASCII 92 (60): '\\'
    rom[1920] = 16'b0000000000000000;
    rom[1921] = 16'b0000000000000000;
    rom[1922] = 16'b0000000000000000;
    rom[1923] = 16'b0000000000000000;
    rom[1924] = 16'b0000000000000000;
    rom[1925] = 16'b0001100000000000;
    rom[1926] = 16'b0000110000000000;
    rom[1927] = 16'b0000110000000000;
    rom[1928] = 16'b0000110000000000;
    rom[1929] = 16'b0000011000000000;
    rom[1930] = 16'b0000011000000000;
    rom[1931] = 16'b0000001100000000;
    rom[1932] = 16'b0000001100000000;
    rom[1933] = 16'b0000001100000000;
    rom[1934] = 16'b0000000110000000;
    rom[1935] = 16'b0000000110000000;
    rom[1936] = 16'b0000000011000000;
    rom[1937] = 16'b0000000011000000;
    rom[1938] = 16'b0000000011000000;
    rom[1939] = 16'b0000000001100000;
    rom[1940] = 16'b0000000001100000;
    rom[1941] = 16'b0000000000110000;
    rom[1942] = 16'b0000000000110000;
    rom[1943] = 16'b0000000000110000;
    rom[1944] = 16'b0000000000011000;
    rom[1945] = 16'b0000000000000000;
    rom[1946] = 16'b0000000000000000;
    rom[1947] = 16'b0000000000000000;
    rom[1948] = 16'b0000000000000000;
    rom[1949] = 16'b0000000000000000;
    rom[1950] = 16'b0000000000000000;
    rom[1951] = 16'b0000000000000000;

    // ASCII 93 (61): ']'
    rom[1952] = 16'b0000000000000000;
    rom[1953] = 16'b0000000000000000;
    rom[1954] = 16'b0000000000000000;
    rom[1955] = 16'b0000000000000000;
    rom[1956] = 16'b0000111111000000;
    rom[1957] = 16'b0000111111000000;
    rom[1958] = 16'b0000000011000000;
    rom[1959] = 16'b0000000011000000;
    rom[1960] = 16'b0000000011000000;
    rom[1961] = 16'b0000000011000000;
    rom[1962] = 16'b0000000011000000;
    rom[1963] = 16'b0000000011000000;
    rom[1964] = 16'b0000000011000000;
    rom[1965] = 16'b0000000011000000;
    rom[1966] = 16'b0000000011000000;
    rom[1967] = 16'b0000000011000000;
    rom[1968] = 16'b0000000011000000;
    rom[1969] = 16'b0000000011000000;
    rom[1970] = 16'b0000000011000000;
    rom[1971] = 16'b0000000011000000;
    rom[1972] = 16'b0000000011000000;
    rom[1973] = 16'b0000000011000000;
    rom[1974] = 16'b0000000011000000;
    rom[1975] = 16'b0000000011000000;
    rom[1976] = 16'b0000111111000000;
    rom[1977] = 16'b0000111111000000;
    rom[1978] = 16'b0000000000000000;
    rom[1979] = 16'b0000000000000000;
    rom[1980] = 16'b0000000000000000;
    rom[1981] = 16'b0000000000000000;
    rom[1982] = 16'b0000000000000000;
    rom[1983] = 16'b0000000000000000;

    // ASCII 94 (62): '^'
    rom[1984] = 16'b0000000000000000;
    rom[1985] = 16'b0000000000000000;
    rom[1986] = 16'b0000000000000000;
    rom[1987] = 16'b0000000000000000;
    rom[1988] = 16'b0000000000000000;
    rom[1989] = 16'b0000000000000000;
    rom[1990] = 16'b0000000000000000;
    rom[1991] = 16'b0000000000000000;
    rom[1992] = 16'b0000000000000000;
    rom[1993] = 16'b0000001110000000;
    rom[1994] = 16'b0000001110000000;
    rom[1995] = 16'b0000011011000000;
    rom[1996] = 16'b0000010001000000;
    rom[1997] = 16'b0000110001100000;
    rom[1998] = 16'b0001100000110000;
    rom[1999] = 16'b0001100000110000;
    rom[2000] = 16'b0000000000000000;
    rom[2001] = 16'b0000000000000000;
    rom[2002] = 16'b0000000000000000;
    rom[2003] = 16'b0000000000000000;
    rom[2004] = 16'b0000000000000000;
    rom[2005] = 16'b0000000000000000;
    rom[2006] = 16'b0000000000000000;
    rom[2007] = 16'b0000000000000000;
    rom[2008] = 16'b0000000000000000;
    rom[2009] = 16'b0000000000000000;
    rom[2010] = 16'b0000000000000000;
    rom[2011] = 16'b0000000000000000;
    rom[2012] = 16'b0000000000000000;
    rom[2013] = 16'b0000000000000000;
    rom[2014] = 16'b0000000000000000;
    rom[2015] = 16'b0000000000000000;

    // ASCII 95 (63): '_'
    rom[2016] = 16'b0000000000000000;
    rom[2017] = 16'b0000000000000000;
    rom[2018] = 16'b0000000000000000;
    rom[2019] = 16'b0000000000000000;
    rom[2020] = 16'b0000000000000000;
    rom[2021] = 16'b0000000000000000;
    rom[2022] = 16'b0000000000000000;
    rom[2023] = 16'b0000000000000000;
    rom[2024] = 16'b0000000000000000;
    rom[2025] = 16'b0000000000000000;
    rom[2026] = 16'b0000000000000000;
    rom[2027] = 16'b0000000000000000;
    rom[2028] = 16'b0000000000000000;
    rom[2029] = 16'b0000000000000000;
    rom[2030] = 16'b0000000000000000;
    rom[2031] = 16'b0000000000000000;
    rom[2032] = 16'b0000000000000000;
    rom[2033] = 16'b0000000000000000;
    rom[2034] = 16'b0000000000000000;
    rom[2035] = 16'b0000000000000000;
    rom[2036] = 16'b0000000000000000;
    rom[2037] = 16'b0000000000000000;
    rom[2038] = 16'b0000000000000000;
    rom[2039] = 16'b0000000000000000;
    rom[2040] = 16'b0000000000000000;
    rom[2041] = 16'b0000000000000000;
    rom[2042] = 16'b0000000000000000;
    rom[2043] = 16'b0000000000000000;
    rom[2044] = 16'b0000000000000000;
    rom[2045] = 16'b0000000000000000;
    rom[2046] = 16'b0000000000000000;
    rom[2047] = 16'b0000000000000000;

    // ASCII 96 (64): '`'
    rom[2048] = 16'b0000000000000000;
    rom[2049] = 16'b0000000000000000;
    rom[2050] = 16'b0000000000000000;
    rom[2051] = 16'b0000000000000000;
    rom[2052] = 16'b0000000000000000;
    rom[2053] = 16'b0000000000000000;
    rom[2054] = 16'b0000111000000000;
    rom[2055] = 16'b0000011100000000;
    rom[2056] = 16'b0000001110000000;
    rom[2057] = 16'b0000000000000000;
    rom[2058] = 16'b0000000000000000;
    rom[2059] = 16'b0000000000000000;
    rom[2060] = 16'b0000000000000000;
    rom[2061] = 16'b0000000000000000;
    rom[2062] = 16'b0000000000000000;
    rom[2063] = 16'b0000000000000000;
    rom[2064] = 16'b0000000000000000;
    rom[2065] = 16'b0000000000000000;
    rom[2066] = 16'b0000000000000000;
    rom[2067] = 16'b0000000000000000;
    rom[2068] = 16'b0000000000000000;
    rom[2069] = 16'b0000000000000000;
    rom[2070] = 16'b0000000000000000;
    rom[2071] = 16'b0000000000000000;
    rom[2072] = 16'b0000000000000000;
    rom[2073] = 16'b0000000000000000;
    rom[2074] = 16'b0000000000000000;
    rom[2075] = 16'b0000000000000000;
    rom[2076] = 16'b0000000000000000;
    rom[2077] = 16'b0000000000000000;
    rom[2078] = 16'b0000000000000000;
    rom[2079] = 16'b0000000000000000;

    // ASCII 97 (65): 'a'
    rom[2080] = 16'b0000000000000000;
    rom[2081] = 16'b0000000000000000;
    rom[2082] = 16'b0000000000000000;
    rom[2083] = 16'b0000000000000000;
    rom[2084] = 16'b0000000000000000;
    rom[2085] = 16'b0000000000000000;
    rom[2086] = 16'b0000000000000000;
    rom[2087] = 16'b0000000000000000;
    rom[2088] = 16'b0000000000000000;
    rom[2089] = 16'b0000000000000000;
    rom[2090] = 16'b0000000000000000;
    rom[2091] = 16'b0000000000000000;
    rom[2092] = 16'b0000000000000000;
    rom[2093] = 16'b0000000000000000;
    rom[2094] = 16'b0000011111100000;
    rom[2095] = 16'b0000111111110000;
    rom[2096] = 16'b0000100000111000;
    rom[2097] = 16'b0000000000011000;
    rom[2098] = 16'b0000000000011000;
    rom[2099] = 16'b0000011111111000;
    rom[2100] = 16'b0000111111111000;
    rom[2101] = 16'b0001110000011000;
    rom[2102] = 16'b0001100000011000;
    rom[2103] = 16'b0001100001111000;
    rom[2104] = 16'b0001111111111000;
    rom[2105] = 16'b0000011110011000;
    rom[2106] = 16'b0000000000000000;
    rom[2107] = 16'b0000000000000000;
    rom[2108] = 16'b0000000000000000;
    rom[2109] = 16'b0000000000000000;
    rom[2110] = 16'b0000000000000000;
    rom[2111] = 16'b0000000000000000;

    // ASCII 98 (66): 'b'
    rom[2112] = 16'b0000000000000000;
    rom[2113] = 16'b0000000000000000;
    rom[2114] = 16'b0000000000000000;
    rom[2115] = 16'b0000000000000000;
    rom[2116] = 16'b0000000000000000;
    rom[2117] = 16'b0000000000000000;
    rom[2118] = 16'b0001100000000000;
    rom[2119] = 16'b0001100000000000;
    rom[2120] = 16'b0001100000000000;
    rom[2121] = 16'b0001100000000000;
    rom[2122] = 16'b0001100000000000;
    rom[2123] = 16'b0001100111100000;
    rom[2124] = 16'b0001111111110000;
    rom[2125] = 16'b0001111000110000;
    rom[2126] = 16'b0001110000011000;
    rom[2127] = 16'b0001100000011000;
    rom[2128] = 16'b0001100000011000;
    rom[2129] = 16'b0001100000011000;
    rom[2130] = 16'b0001100000011000;
    rom[2131] = 16'b0001100000111000;
    rom[2132] = 16'b0001100001110000;
    rom[2133] = 16'b0001111111100000;
    rom[2134] = 16'b0000111111000000;
    rom[2135] = 16'b0000000000000000;
    rom[2136] = 16'b0000000000000000;
    rom[2137] = 16'b0000000000000000;
    rom[2138] = 16'b0000000000000000;
    rom[2139] = 16'b0000000000000000;
    rom[2140] = 16'b0000000000000000;
    rom[2141] = 16'b0000000000000000;
    rom[2142] = 16'b0000000000000000;
    rom[2143] = 16'b0000000000000000;

    // ASCII 99 (67): 'c'
    rom[2144] = 16'b0000000000000000;
    rom[2145] = 16'b0000000000000000;
    rom[2146] = 16'b0000000000000000;
    rom[2147] = 16'b0000000000000000;
    rom[2148] = 16'b0000000000000000;
    rom[2149] = 16'b0000000000000000;
    rom[2150] = 16'b0000000000000000;
    rom[2151] = 16'b0000000000000000;
    rom[2152] = 16'b0000000000000000;
    rom[2153] = 16'b0000000000000000;
    rom[2154] = 16'b0000000000000000;
    rom[2155] = 16'b0000000000000000;
    rom[2156] = 16'b0000000000000000;
    rom[2157] = 16'b0000000000000000;
    rom[2158] = 16'b0000001111100000;
    rom[2159] = 16'b0000011111110000;
    rom[2160] = 16'b0000111000010000;
    rom[2161] = 16'b0001110000000000;
    rom[2162] = 16'b0001100000000000;
    rom[2163] = 16'b0001100000000000;
    rom[2164] = 16'b0001100000000000;
    rom[2165] = 16'b0001100000000000;
    rom[2166] = 16'b0001110000000000;
    rom[2167] = 16'b0000111000010000;
    rom[2168] = 16'b0000111111110000;
    rom[2169] = 16'b0000001111100000;
    rom[2170] = 16'b0000000000000000;
    rom[2171] = 16'b0000000000000000;
    rom[2172] = 16'b0000000000000000;
    rom[2173] = 16'b0000000000000000;
    rom[2174] = 16'b0000000000000000;
    rom[2175] = 16'b0000000000000000;

    // ASCII 100 (68): 'd'
    rom[2176] = 16'b0000000000000000;
    rom[2177] = 16'b0000000000000000;
    rom[2178] = 16'b0000000000000000;
    rom[2179] = 16'b0000000000000000;
    rom[2180] = 16'b0000000000000000;
    rom[2181] = 16'b0000000000000000;
    rom[2182] = 16'b0000000000110000;
    rom[2183] = 16'b0000000000110000;
    rom[2184] = 16'b0000000000110000;
    rom[2185] = 16'b0000000000110000;
    rom[2186] = 16'b0000000000110000;
    rom[2187] = 16'b0000011111110000;
    rom[2188] = 16'b0000111111110000;
    rom[2189] = 16'b0001110000110000;
    rom[2190] = 16'b0011100000110000;
    rom[2191] = 16'b0011000000110000;
    rom[2192] = 16'b0011000000110000;
    rom[2193] = 16'b0011000000110000;
    rom[2194] = 16'b0011000000110000;
    rom[2195] = 16'b0011000001110000;
    rom[2196] = 16'b0001100011110000;
    rom[2197] = 16'b0001111110110000;
    rom[2198] = 16'b0000111100110000;
    rom[2199] = 16'b0000000000000000;
    rom[2200] = 16'b0000000000000000;
    rom[2201] = 16'b0000000000000000;
    rom[2202] = 16'b0000000000000000;
    rom[2203] = 16'b0000000000000000;
    rom[2204] = 16'b0000000000000000;
    rom[2205] = 16'b0000000000000000;
    rom[2206] = 16'b0000000000000000;
    rom[2207] = 16'b0000000000000000;

    // ASCII 101 (69): 'e'
    rom[2208] = 16'b0000000000000000;
    rom[2209] = 16'b0000000000000000;
    rom[2210] = 16'b0000000000000000;
    rom[2211] = 16'b0000000000000000;
    rom[2212] = 16'b0000000000000000;
    rom[2213] = 16'b0000000000000000;
    rom[2214] = 16'b0000000000000000;
    rom[2215] = 16'b0000000000000000;
    rom[2216] = 16'b0000000000000000;
    rom[2217] = 16'b0000000000000000;
    rom[2218] = 16'b0000000000000000;
    rom[2219] = 16'b0000000000000000;
    rom[2220] = 16'b0000000000000000;
    rom[2221] = 16'b0000000000000000;
    rom[2222] = 16'b0000011110000000;
    rom[2223] = 16'b0000111111100000;
    rom[2224] = 16'b0001100001100000;
    rom[2225] = 16'b0011000000110000;
    rom[2226] = 16'b0011000000110000;
    rom[2227] = 16'b0011111111110000;
    rom[2228] = 16'b0011111111110000;
    rom[2229] = 16'b0011000000000000;
    rom[2230] = 16'b0011000000000000;
    rom[2231] = 16'b0001100000100000;
    rom[2232] = 16'b0001111111100000;
    rom[2233] = 16'b0000011111000000;
    rom[2234] = 16'b0000000000000000;
    rom[2235] = 16'b0000000000000000;
    rom[2236] = 16'b0000000000000000;
    rom[2237] = 16'b0000000000000000;
    rom[2238] = 16'b0000000000000000;
    rom[2239] = 16'b0000000000000000;

    // ASCII 102 (70): 'f'
    rom[2240] = 16'b0000000000000000;
    rom[2241] = 16'b0000000000000000;
    rom[2242] = 16'b0000000000000000;
    rom[2243] = 16'b0000000000000000;
    rom[2244] = 16'b0000000000000000;
    rom[2245] = 16'b0000000000000000;
    rom[2246] = 16'b0000000011111000;
    rom[2247] = 16'b0000000111111000;
    rom[2248] = 16'b0000001110000000;
    rom[2249] = 16'b0000001100000000;
    rom[2250] = 16'b0000001100000000;
    rom[2251] = 16'b0000001100000000;
    rom[2252] = 16'b0011111111110000;
    rom[2253] = 16'b0011111111110000;
    rom[2254] = 16'b0000001100000000;
    rom[2255] = 16'b0000001100000000;
    rom[2256] = 16'b0000001100000000;
    rom[2257] = 16'b0000001100000000;
    rom[2258] = 16'b0000001100000000;
    rom[2259] = 16'b0000001100000000;
    rom[2260] = 16'b0000001100000000;
    rom[2261] = 16'b0000001100000000;
    rom[2262] = 16'b0000001100000000;
    rom[2263] = 16'b0000000000000000;
    rom[2264] = 16'b0000000000000000;
    rom[2265] = 16'b0000000000000000;
    rom[2266] = 16'b0000000000000000;
    rom[2267] = 16'b0000000000000000;
    rom[2268] = 16'b0000000000000000;
    rom[2269] = 16'b0000000000000000;
    rom[2270] = 16'b0000000000000000;
    rom[2271] = 16'b0000000000000000;

    // ASCII 103 (71): 'g'
    rom[2272] = 16'b0000000000000000;
    rom[2273] = 16'b0000000000000000;
    rom[2274] = 16'b0000000000000000;
    rom[2275] = 16'b0000000000000000;
    rom[2276] = 16'b0000000000000000;
    rom[2277] = 16'b0000000000000000;
    rom[2278] = 16'b0000000000000000;
    rom[2279] = 16'b0000000000000000;
    rom[2280] = 16'b0000000000000000;
    rom[2281] = 16'b0000000000000000;
    rom[2282] = 16'b0000000000000000;
    rom[2283] = 16'b0000011111111000;
    rom[2284] = 16'b0000111111111000;
    rom[2285] = 16'b0001110001110000;
    rom[2286] = 16'b0001100000110000;
    rom[2287] = 16'b0001100000110000;
    rom[2288] = 16'b0001110001110000;
    rom[2289] = 16'b0000111111100000;
    rom[2290] = 16'b0001111111000000;
    rom[2291] = 16'b0011000000000000;
    rom[2292] = 16'b0011000000000000;
    rom[2293] = 16'b0001111111100000;
    rom[2294] = 16'b0001111111111000;
    rom[2295] = 16'b0011000000011000;
    rom[2296] = 16'b0011000000011000;
    rom[2297] = 16'b0011100000111000;
    rom[2298] = 16'b0011111111110000;
    rom[2299] = 16'b0000111111000000;
    rom[2300] = 16'b0000000000000000;
    rom[2301] = 16'b0000000000000000;
    rom[2302] = 16'b0000000000000000;
    rom[2303] = 16'b0000000000000000;

    // ASCII 104 (72): 'h'
    rom[2304] = 16'b0000000000000000;
    rom[2305] = 16'b0000000000000000;
    rom[2306] = 16'b0000000000000000;
    rom[2307] = 16'b0000000000000000;
    rom[2308] = 16'b0000000000000000;
    rom[2309] = 16'b0000000000000000;
    rom[2310] = 16'b0001100000000000;
    rom[2311] = 16'b0001100000000000;
    rom[2312] = 16'b0001100000000000;
    rom[2313] = 16'b0001100000000000;
    rom[2314] = 16'b0001100000000000;
    rom[2315] = 16'b0001100111000000;
    rom[2316] = 16'b0001111111100000;
    rom[2317] = 16'b0001111001110000;
    rom[2318] = 16'b0001110000110000;
    rom[2319] = 16'b0001100000110000;
    rom[2320] = 16'b0001100000110000;
    rom[2321] = 16'b0001100000110000;
    rom[2322] = 16'b0001100000110000;
    rom[2323] = 16'b0001100000110000;
    rom[2324] = 16'b0001100000110000;
    rom[2325] = 16'b0001100000110000;
    rom[2326] = 16'b0001100000110000;
    rom[2327] = 16'b0000000000000000;
    rom[2328] = 16'b0000000000000000;
    rom[2329] = 16'b0000000000000000;
    rom[2330] = 16'b0000000000000000;
    rom[2331] = 16'b0000000000000000;
    rom[2332] = 16'b0000000000000000;
    rom[2333] = 16'b0000000000000000;
    rom[2334] = 16'b0000000000000000;
    rom[2335] = 16'b0000000000000000;

    // ASCII 105 (73): 'i'
    rom[2336] = 16'b0000000000000000;
    rom[2337] = 16'b0000000000000000;
    rom[2338] = 16'b0000000000000000;
    rom[2339] = 16'b0000000000000000;
    rom[2340] = 16'b0000000000000000;
    rom[2341] = 16'b0000000000000000;
    rom[2342] = 16'b0000001110000000;
    rom[2343] = 16'b0000001110000000;
    rom[2344] = 16'b0000001110000000;
    rom[2345] = 16'b0000000000000000;
    rom[2346] = 16'b0000000000000000;
    rom[2347] = 16'b0001111110000000;
    rom[2348] = 16'b0001111110000000;
    rom[2349] = 16'b0000000110000000;
    rom[2350] = 16'b0000000110000000;
    rom[2351] = 16'b0000000110000000;
    rom[2352] = 16'b0000000110000000;
    rom[2353] = 16'b0000000110000000;
    rom[2354] = 16'b0000000110000000;
    rom[2355] = 16'b0000000110000000;
    rom[2356] = 16'b0000000110000000;
    rom[2357] = 16'b0001111111110000;
    rom[2358] = 16'b0001111111110000;
    rom[2359] = 16'b0000000000000000;
    rom[2360] = 16'b0000000000000000;
    rom[2361] = 16'b0000000000000000;
    rom[2362] = 16'b0000000000000000;
    rom[2363] = 16'b0000000000000000;
    rom[2364] = 16'b0000000000000000;
    rom[2365] = 16'b0000000000000000;
    rom[2366] = 16'b0000000000000000;
    rom[2367] = 16'b0000000000000000;

    // ASCII 106 (74): 'j'
    rom[2368] = 16'b0000000000000000;
    rom[2369] = 16'b0000000000000000;
    rom[2370] = 16'b0000000000000000;
    rom[2371] = 16'b0000000000000000;
    rom[2372] = 16'b0000000011100000;
    rom[2373] = 16'b0000000011100000;
    rom[2374] = 16'b0000000011100000;
    rom[2375] = 16'b0000000000000000;
    rom[2376] = 16'b0000000000000000;
    rom[2377] = 16'b0001111111100000;
    rom[2378] = 16'b0001111111100000;
    rom[2379] = 16'b0000000001100000;
    rom[2380] = 16'b0000000001100000;
    rom[2381] = 16'b0000000001100000;
    rom[2382] = 16'b0000000001100000;
    rom[2383] = 16'b0000000001100000;
    rom[2384] = 16'b0000000001100000;
    rom[2385] = 16'b0000000001100000;
    rom[2386] = 16'b0000000001100000;
    rom[2387] = 16'b0000000001100000;
    rom[2388] = 16'b0000000001100000;
    rom[2389] = 16'b0000000001100000;
    rom[2390] = 16'b0000000001100000;
    rom[2391] = 16'b0001000011000000;
    rom[2392] = 16'b0001111111000000;
    rom[2393] = 16'b0000111100000000;
    rom[2394] = 16'b0000000000000000;
    rom[2395] = 16'b0000000000000000;
    rom[2396] = 16'b0000000000000000;
    rom[2397] = 16'b0000000000000000;
    rom[2398] = 16'b0000000000000000;
    rom[2399] = 16'b0000000000000000;

    // ASCII 107 (75): 'k'
    rom[2400] = 16'b0000000000000000;
    rom[2401] = 16'b0000000000000000;
    rom[2402] = 16'b0000000000000000;
    rom[2403] = 16'b0000000000000000;
    rom[2404] = 16'b0000000000000000;
    rom[2405] = 16'b0000000000000000;
    rom[2406] = 16'b0001100000000000;
    rom[2407] = 16'b0001100000000000;
    rom[2408] = 16'b0001100000000000;
    rom[2409] = 16'b0001100000000000;
    rom[2410] = 16'b0001100000000000;
    rom[2411] = 16'b0001100000111000;
    rom[2412] = 16'b0001100001110000;
    rom[2413] = 16'b0001100011100000;
    rom[2414] = 16'b0001100111000000;
    rom[2415] = 16'b0001101100000000;
    rom[2416] = 16'b0001111000000000;
    rom[2417] = 16'b0001101100000000;
    rom[2418] = 16'b0001100110000000;
    rom[2419] = 16'b0001100011000000;
    rom[2420] = 16'b0001100001100000;
    rom[2421] = 16'b0001100000110000;
    rom[2422] = 16'b0001100000011000;
    rom[2423] = 16'b0000000000000000;
    rom[2424] = 16'b0000000000000000;
    rom[2425] = 16'b0000000000000000;
    rom[2426] = 16'b0000000000000000;
    rom[2427] = 16'b0000000000000000;
    rom[2428] = 16'b0000000000000000;
    rom[2429] = 16'b0000000000000000;
    rom[2430] = 16'b0000000000000000;
    rom[2431] = 16'b0000000000000000;

    // ASCII 108 (76): 'l'
    rom[2432] = 16'b0000000000000000;
    rom[2433] = 16'b0000000000000000;
    rom[2434] = 16'b0000000000000000;
    rom[2435] = 16'b0000000000000000;
    rom[2436] = 16'b0000000000000000;
    rom[2437] = 16'b0000000000000000;
    rom[2438] = 16'b0001111110000000;
    rom[2439] = 16'b0001111110000000;
    rom[2440] = 16'b0000000110000000;
    rom[2441] = 16'b0000000110000000;
    rom[2442] = 16'b0000000110000000;
    rom[2443] = 16'b0000000110000000;
    rom[2444] = 16'b0000000110000000;
    rom[2445] = 16'b0000000110000000;
    rom[2446] = 16'b0000000110000000;
    rom[2447] = 16'b0000000110000000;
    rom[2448] = 16'b0000000110000000;
    rom[2449] = 16'b0000000110000000;
    rom[2450] = 16'b0000000110000000;
    rom[2451] = 16'b0000000110000000;
    rom[2452] = 16'b0000000110000000;
    rom[2453] = 16'b0001111111110000;
    rom[2454] = 16'b0001111111110000;
    rom[2455] = 16'b0000000000000000;
    rom[2456] = 16'b0000000000000000;
    rom[2457] = 16'b0000000000000000;
    rom[2458] = 16'b0000000000000000;
    rom[2459] = 16'b0000000000000000;
    rom[2460] = 16'b0000000000000000;
    rom[2461] = 16'b0000000000000000;
    rom[2462] = 16'b0000000000000000;
    rom[2463] = 16'b0000000000000000;

    // ASCII 109 (77): 'm'
    rom[2464] = 16'b0000000000000000;
    rom[2465] = 16'b0000000000000000;
    rom[2466] = 16'b0000000000000000;
    rom[2467] = 16'b0000000000000000;
    rom[2468] = 16'b0000000000000000;
    rom[2469] = 16'b0000000000000000;
    rom[2470] = 16'b0000000000000000;
    rom[2471] = 16'b0000000000000000;
    rom[2472] = 16'b0000000000000000;
    rom[2473] = 16'b0000000000000000;
    rom[2474] = 16'b0000000000000000;
    rom[2475] = 16'b0000000000000000;
    rom[2476] = 16'b0000000000000000;
    rom[2477] = 16'b0000000000000000;
    rom[2478] = 16'b0011011100111000;
    rom[2479] = 16'b0011111111111100;
    rom[2480] = 16'b0011100111001100;
    rom[2481] = 16'b0011100111001100;
    rom[2482] = 16'b0011000110001100;
    rom[2483] = 16'b0011000110001100;
    rom[2484] = 16'b0011000110001100;
    rom[2485] = 16'b0011000110001100;
    rom[2486] = 16'b0011000110001100;
    rom[2487] = 16'b0011000110001100;
    rom[2488] = 16'b0011000110001100;
    rom[2489] = 16'b0011000110001100;
    rom[2490] = 16'b0000000000000000;
    rom[2491] = 16'b0000000000000000;
    rom[2492] = 16'b0000000000000000;
    rom[2493] = 16'b0000000000000000;
    rom[2494] = 16'b0000000000000000;
    rom[2495] = 16'b0000000000000000;

    // ASCII 110 (78): 'n'
    rom[2496] = 16'b0000000000000000;
    rom[2497] = 16'b0000000000000000;
    rom[2498] = 16'b0000000000000000;
    rom[2499] = 16'b0000000000000000;
    rom[2500] = 16'b0000000000000000;
    rom[2501] = 16'b0000000000000000;
    rom[2502] = 16'b0000000000000000;
    rom[2503] = 16'b0000000000000000;
    rom[2504] = 16'b0000000000000000;
    rom[2505] = 16'b0000000000000000;
    rom[2506] = 16'b0000000000000000;
    rom[2507] = 16'b0000000000000000;
    rom[2508] = 16'b0000000000000000;
    rom[2509] = 16'b0000000000000000;
    rom[2510] = 16'b0001100111000000;
    rom[2511] = 16'b0001111111100000;
    rom[2512] = 16'b0001111001110000;
    rom[2513] = 16'b0001110000110000;
    rom[2514] = 16'b0001100000110000;
    rom[2515] = 16'b0001100000110000;
    rom[2516] = 16'b0001100000110000;
    rom[2517] = 16'b0001100000110000;
    rom[2518] = 16'b0001100000110000;
    rom[2519] = 16'b0001100000110000;
    rom[2520] = 16'b0001100000110000;
    rom[2521] = 16'b0001100000110000;
    rom[2522] = 16'b0000000000000000;
    rom[2523] = 16'b0000000000000000;
    rom[2524] = 16'b0000000000000000;
    rom[2525] = 16'b0000000000000000;
    rom[2526] = 16'b0000000000000000;
    rom[2527] = 16'b0000000000000000;

    // ASCII 111 (79): 'o'
    rom[2528] = 16'b0000000000000000;
    rom[2529] = 16'b0000000000000000;
    rom[2530] = 16'b0000000000000000;
    rom[2531] = 16'b0000000000000000;
    rom[2532] = 16'b0000000000000000;
    rom[2533] = 16'b0000000000000000;
    rom[2534] = 16'b0000000000000000;
    rom[2535] = 16'b0000000000000000;
    rom[2536] = 16'b0000000000000000;
    rom[2537] = 16'b0000000000000000;
    rom[2538] = 16'b0000000000000000;
    rom[2539] = 16'b0000000000000000;
    rom[2540] = 16'b0000000000000000;
    rom[2541] = 16'b0000000000000000;
    rom[2542] = 16'b0000011111000000;
    rom[2543] = 16'b0000111111110000;
    rom[2544] = 16'b0001110001110000;
    rom[2545] = 16'b0011100000111000;
    rom[2546] = 16'b0011000000011000;
    rom[2547] = 16'b0011000000011000;
    rom[2548] = 16'b0011000000011000;
    rom[2549] = 16'b0011000000011000;
    rom[2550] = 16'b0011100000111000;
    rom[2551] = 16'b0001110001110000;
    rom[2552] = 16'b0001111111100000;
    rom[2553] = 16'b0000011111000000;
    rom[2554] = 16'b0000000000000000;
    rom[2555] = 16'b0000000000000000;
    rom[2556] = 16'b0000000000000000;
    rom[2557] = 16'b0000000000000000;
    rom[2558] = 16'b0000000000000000;
    rom[2559] = 16'b0000000000000000;

    // ASCII 112 (80): 'p'
    rom[2560] = 16'b0000000000000000;
    rom[2561] = 16'b0000000000000000;
    rom[2562] = 16'b0000000000000000;
    rom[2563] = 16'b0000000000000000;
    rom[2564] = 16'b0000000000000000;
    rom[2565] = 16'b0000000000000000;
    rom[2566] = 16'b0000000000000000;
    rom[2567] = 16'b0000000000000000;
    rom[2568] = 16'b0000000000000000;
    rom[2569] = 16'b0000000000000000;
    rom[2570] = 16'b0000000000000000;
    rom[2571] = 16'b0001100111100000;
    rom[2572] = 16'b0001111111110000;
    rom[2573] = 16'b0001111000110000;
    rom[2574] = 16'b0001110000011000;
    rom[2575] = 16'b0001100000011000;
    rom[2576] = 16'b0001100000011000;
    rom[2577] = 16'b0001100000011000;
    rom[2578] = 16'b0001100000011000;
    rom[2579] = 16'b0001100000111000;
    rom[2580] = 16'b0001100001110000;
    rom[2581] = 16'b0001111111100000;
    rom[2582] = 16'b0001111111000000;
    rom[2583] = 16'b0001100000000000;
    rom[2584] = 16'b0001100000000000;
    rom[2585] = 16'b0001100000000000;
    rom[2586] = 16'b0001100000000000;
    rom[2587] = 16'b0001100000000000;
    rom[2588] = 16'b0000000000000000;
    rom[2589] = 16'b0000000000000000;
    rom[2590] = 16'b0000000000000000;
    rom[2591] = 16'b0000000000000000;

    // ASCII 113 (81): 'q'
    rom[2592] = 16'b0000000000000000;
    rom[2593] = 16'b0000000000000000;
    rom[2594] = 16'b0000000000000000;
    rom[2595] = 16'b0000000000000000;
    rom[2596] = 16'b0000000000000000;
    rom[2597] = 16'b0000000000000000;
    rom[2598] = 16'b0000000000000000;
    rom[2599] = 16'b0000000000000000;
    rom[2600] = 16'b0000000000000000;
    rom[2601] = 16'b0000000000000000;
    rom[2602] = 16'b0000000000000000;
    rom[2603] = 16'b0000011111110000;
    rom[2604] = 16'b0000111111110000;
    rom[2605] = 16'b0001110000110000;
    rom[2606] = 16'b0011100000110000;
    rom[2607] = 16'b0011000000110000;
    rom[2608] = 16'b0011000000110000;
    rom[2609] = 16'b0011000000110000;
    rom[2610] = 16'b0011000000110000;
    rom[2611] = 16'b0011000001110000;
    rom[2612] = 16'b0001100011110000;
    rom[2613] = 16'b0001111110110000;
    rom[2614] = 16'b0000111100110000;
    rom[2615] = 16'b0000000000110000;
    rom[2616] = 16'b0000000000110000;
    rom[2617] = 16'b0000000000110000;
    rom[2618] = 16'b0000000000110000;
    rom[2619] = 16'b0000000000110000;
    rom[2620] = 16'b0000000000000000;
    rom[2621] = 16'b0000000000000000;
    rom[2622] = 16'b0000000000000000;
    rom[2623] = 16'b0000000000000000;

    // ASCII 114 (82): 'r'
    rom[2624] = 16'b0000000000000000;
    rom[2625] = 16'b0000000000000000;
    rom[2626] = 16'b0000000000000000;
    rom[2627] = 16'b0000000000000000;
    rom[2628] = 16'b0000000000000000;
    rom[2629] = 16'b0000000000000000;
    rom[2630] = 16'b0000000000000000;
    rom[2631] = 16'b0000000000000000;
    rom[2632] = 16'b0000000000000000;
    rom[2633] = 16'b0000000000000000;
    rom[2634] = 16'b0000000000000000;
    rom[2635] = 16'b0000000000000000;
    rom[2636] = 16'b0000000000000000;
    rom[2637] = 16'b0000000000000000;
    rom[2638] = 16'b0001100111100000;
    rom[2639] = 16'b0001101111110000;
    rom[2640] = 16'b0001111000111000;
    rom[2641] = 16'b0001110000011000;
    rom[2642] = 16'b0001100000011000;
    rom[2643] = 16'b0001100000000000;
    rom[2644] = 16'b0001100000000000;
    rom[2645] = 16'b0001100000000000;
    rom[2646] = 16'b0001100000000000;
    rom[2647] = 16'b0001100000000000;
    rom[2648] = 16'b0001100000000000;
    rom[2649] = 16'b0001100000000000;
    rom[2650] = 16'b0000000000000000;
    rom[2651] = 16'b0000000000000000;
    rom[2652] = 16'b0000000000000000;
    rom[2653] = 16'b0000000000000000;
    rom[2654] = 16'b0000000000000000;
    rom[2655] = 16'b0000000000000000;

    // ASCII 115 (83): 's'
    rom[2656] = 16'b0000000000000000;
    rom[2657] = 16'b0000000000000000;
    rom[2658] = 16'b0000000000000000;
    rom[2659] = 16'b0000000000000000;
    rom[2660] = 16'b0000000000000000;
    rom[2661] = 16'b0000000000000000;
    rom[2662] = 16'b0000000000000000;
    rom[2663] = 16'b0000000000000000;
    rom[2664] = 16'b0000000000000000;
    rom[2665] = 16'b0000000000000000;
    rom[2666] = 16'b0000000000000000;
    rom[2667] = 16'b0000000000000000;
    rom[2668] = 16'b0000000000000000;
    rom[2669] = 16'b0000000000000000;
    rom[2670] = 16'b0000011111000000;
    rom[2671] = 16'b0000111111100000;
    rom[2672] = 16'b0001100000100000;
    rom[2673] = 16'b0001100000000000;
    rom[2674] = 16'b0001110000000000;
    rom[2675] = 16'b0000111110000000;
    rom[2676] = 16'b0000001111100000;
    rom[2677] = 16'b0000000001110000;
    rom[2678] = 16'b0000000000110000;
    rom[2679] = 16'b0001000000110000;
    rom[2680] = 16'b0001111111100000;
    rom[2681] = 16'b0000111111000000;
    rom[2682] = 16'b0000000000000000;
    rom[2683] = 16'b0000000000000000;
    rom[2684] = 16'b0000000000000000;
    rom[2685] = 16'b0000000000000000;
    rom[2686] = 16'b0000000000000000;
    rom[2687] = 16'b0000000000000000;

    // ASCII 116 (84): 't'
    rom[2688] = 16'b0000000000000000;
    rom[2689] = 16'b0000000000000000;
    rom[2690] = 16'b0000000000000000;
    rom[2691] = 16'b0000000000000000;
    rom[2692] = 16'b0000000000000000;
    rom[2693] = 16'b0000000000000000;
    rom[2694] = 16'b0000000000000000;
    rom[2695] = 16'b0000000000000000;
    rom[2696] = 16'b0000001000000000;
    rom[2697] = 16'b0000011000000000;
    rom[2698] = 16'b0000011000000000;
    rom[2699] = 16'b0000011000000000;
    rom[2700] = 16'b0011111111111000;
    rom[2701] = 16'b0011111111111000;
    rom[2702] = 16'b0000011000000000;
    rom[2703] = 16'b0000011000000000;
    rom[2704] = 16'b0000011000000000;
    rom[2705] = 16'b0000011000000000;
    rom[2706] = 16'b0000011000000000;
    rom[2707] = 16'b0000011000000000;
    rom[2708] = 16'b0000011100000000;
    rom[2709] = 16'b0000001100000000;
    rom[2710] = 16'b0000001111111000;
    rom[2711] = 16'b0000000111111000;
    rom[2712] = 16'b0000000000000000;
    rom[2713] = 16'b0000000000000000;
    rom[2714] = 16'b0000000000000000;
    rom[2715] = 16'b0000000000000000;
    rom[2716] = 16'b0000000000000000;
    rom[2717] = 16'b0000000000000000;
    rom[2718] = 16'b0000000000000000;
    rom[2719] = 16'b0000000000000000;

    // ASCII 117 (85): 'u'
    rom[2720] = 16'b0000000000000000;
    rom[2721] = 16'b0000000000000000;
    rom[2722] = 16'b0000000000000000;
    rom[2723] = 16'b0000000000000000;
    rom[2724] = 16'b0000000000000000;
    rom[2725] = 16'b0000000000000000;
    rom[2726] = 16'b0000000000000000;
    rom[2727] = 16'b0000000000000000;
    rom[2728] = 16'b0000000000000000;
    rom[2729] = 16'b0000000000000000;
    rom[2730] = 16'b0000000000000000;
    rom[2731] = 16'b0000000000000000;
    rom[2732] = 16'b0000000000000000;
    rom[2733] = 16'b0000000000000000;
    rom[2734] = 16'b0001100000110000;
    rom[2735] = 16'b0001100000110000;
    rom[2736] = 16'b0001100000110000;
    rom[2737] = 16'b0001100000110000;
    rom[2738] = 16'b0001100000110000;
    rom[2739] = 16'b0001100000110000;
    rom[2740] = 16'b0001100000110000;
    rom[2741] = 16'b0001100000110000;
    rom[2742] = 16'b0001100001110000;
    rom[2743] = 16'b0001110011110000;
    rom[2744] = 16'b0000111111110000;
    rom[2745] = 16'b0000111100110000;
    rom[2746] = 16'b0000000000000000;
    rom[2747] = 16'b0000000000000000;
    rom[2748] = 16'b0000000000000000;
    rom[2749] = 16'b0000000000000000;
    rom[2750] = 16'b0000000000000000;
    rom[2751] = 16'b0000000000000000;

    // ASCII 118 (86): 'v'
    rom[2752] = 16'b0000000000000000;
    rom[2753] = 16'b0000000000000000;
    rom[2754] = 16'b0000000000000000;
    rom[2755] = 16'b0000000000000000;
    rom[2756] = 16'b0000000000000000;
    rom[2757] = 16'b0000000000000000;
    rom[2758] = 16'b0000000000000000;
    rom[2759] = 16'b0000000000000000;
    rom[2760] = 16'b0000000000000000;
    rom[2761] = 16'b0000000000000000;
    rom[2762] = 16'b0000000000000000;
    rom[2763] = 16'b0000000000000000;
    rom[2764] = 16'b0000000000000000;
    rom[2765] = 16'b0000000000000000;
    rom[2766] = 16'b0011000000011000;
    rom[2767] = 16'b0011000000011000;
    rom[2768] = 16'b0011100000110000;
    rom[2769] = 16'b0001100000110000;
    rom[2770] = 16'b0001100000110000;
    rom[2771] = 16'b0000110001100000;
    rom[2772] = 16'b0000110001100000;
    rom[2773] = 16'b0000110001000000;
    rom[2774] = 16'b0000011011000000;
    rom[2775] = 16'b0000011011000000;
    rom[2776] = 16'b0000001010000000;
    rom[2777] = 16'b0000001110000000;
    rom[2778] = 16'b0000000000000000;
    rom[2779] = 16'b0000000000000000;
    rom[2780] = 16'b0000000000000000;
    rom[2781] = 16'b0000000000000000;
    rom[2782] = 16'b0000000000000000;
    rom[2783] = 16'b0000000000000000;

    // ASCII 119 (87): 'w'
    rom[2784] = 16'b0000000000000000;
    rom[2785] = 16'b0000000000000000;
    rom[2786] = 16'b0000000000000000;
    rom[2787] = 16'b0000000000000000;
    rom[2788] = 16'b0000000000000000;
    rom[2789] = 16'b0000000000000000;
    rom[2790] = 16'b0000000000000000;
    rom[2791] = 16'b0000000000000000;
    rom[2792] = 16'b0000000000000000;
    rom[2793] = 16'b0000000000000000;
    rom[2794] = 16'b0000000000000000;
    rom[2795] = 16'b0000000000000000;
    rom[2796] = 16'b0000000000000000;
    rom[2797] = 16'b0000000000000000;
    rom[2798] = 16'b0011000000011000;
    rom[2799] = 16'b0011000000011000;
    rom[2800] = 16'b0011000000011000;
    rom[2801] = 16'b0011000100011000;
    rom[2802] = 16'b0011001110011000;
    rom[2803] = 16'b0011001010011000;
    rom[2804] = 16'b0011001010011000;
    rom[2805] = 16'b0011011011011000;
    rom[2806] = 16'b0001011011010000;
    rom[2807] = 16'b0001010001010000;
    rom[2808] = 16'b0001110001110000;
    rom[2809] = 16'b0001110001110000;
    rom[2810] = 16'b0000000000000000;
    rom[2811] = 16'b0000000000000000;
    rom[2812] = 16'b0000000000000000;
    rom[2813] = 16'b0000000000000000;
    rom[2814] = 16'b0000000000000000;
    rom[2815] = 16'b0000000000000000;

    // ASCII 120 (88): 'x'
    rom[2816] = 16'b0000000000000000;
    rom[2817] = 16'b0000000000000000;
    rom[2818] = 16'b0000000000000000;
    rom[2819] = 16'b0000000000000000;
    rom[2820] = 16'b0000000000000000;
    rom[2821] = 16'b0000000000000000;
    rom[2822] = 16'b0000000000000000;
    rom[2823] = 16'b0000000000000000;
    rom[2824] = 16'b0000000000000000;
    rom[2825] = 16'b0000000000000000;
    rom[2826] = 16'b0000000000000000;
    rom[2827] = 16'b0000000000000000;
    rom[2828] = 16'b0000000000000000;
    rom[2829] = 16'b0000000000000000;
    rom[2830] = 16'b0011100000111000;
    rom[2831] = 16'b0001110001110000;
    rom[2832] = 16'b0000110001100000;
    rom[2833] = 16'b0000111011100000;
    rom[2834] = 16'b0000011111000000;
    rom[2835] = 16'b0000001110000000;
    rom[2836] = 16'b0000001110000000;
    rom[2837] = 16'b0000011011000000;
    rom[2838] = 16'b0000111011100000;
    rom[2839] = 16'b0000110001100000;
    rom[2840] = 16'b0001110001110000;
    rom[2841] = 16'b0011100000111000;
    rom[2842] = 16'b0000000000000000;
    rom[2843] = 16'b0000000000000000;
    rom[2844] = 16'b0000000000000000;
    rom[2845] = 16'b0000000000000000;
    rom[2846] = 16'b0000000000000000;
    rom[2847] = 16'b0000000000000000;

    // ASCII 121 (89): 'y'
    rom[2848] = 16'b0000000000000000;
    rom[2849] = 16'b0000000000000000;
    rom[2850] = 16'b0000000000000000;
    rom[2851] = 16'b0000000000000000;
    rom[2852] = 16'b0000000000000000;
    rom[2853] = 16'b0000000000000000;
    rom[2854] = 16'b0000000000000000;
    rom[2855] = 16'b0000000000000000;
    rom[2856] = 16'b0000000000000000;
    rom[2857] = 16'b0000000000000000;
    rom[2858] = 16'b0000000000000000;
    rom[2859] = 16'b0011000000011000;
    rom[2860] = 16'b0011000000011000;
    rom[2861] = 16'b0011100000110000;
    rom[2862] = 16'b0001100000110000;
    rom[2863] = 16'b0001100000110000;
    rom[2864] = 16'b0000110001100000;
    rom[2865] = 16'b0000110001100000;
    rom[2866] = 16'b0000111011000000;
    rom[2867] = 16'b0000011011000000;
    rom[2868] = 16'b0000011010000000;
    rom[2869] = 16'b0000001110000000;
    rom[2870] = 16'b0000001110000000;
    rom[2871] = 16'b0000001100000000;
    rom[2872] = 16'b0000011100000000;
    rom[2873] = 16'b0000111000000000;
    rom[2874] = 16'b0111110000000000;
    rom[2875] = 16'b0111100000000000;
    rom[2876] = 16'b0000000000000000;
    rom[2877] = 16'b0000000000000000;
    rom[2878] = 16'b0000000000000000;
    rom[2879] = 16'b0000000000000000;

    // ASCII 122 (90): 'z'
    rom[2880] = 16'b0000000000000000;
    rom[2881] = 16'b0000000000000000;
    rom[2882] = 16'b0000000000000000;
    rom[2883] = 16'b0000000000000000;
    rom[2884] = 16'b0000000000000000;
    rom[2885] = 16'b0000000000000000;
    rom[2886] = 16'b0000000000000000;
    rom[2887] = 16'b0000000000000000;
    rom[2888] = 16'b0000000000000000;
    rom[2889] = 16'b0000000000000000;
    rom[2890] = 16'b0000000000000000;
    rom[2891] = 16'b0000000000000000;
    rom[2892] = 16'b0000000000000000;
    rom[2893] = 16'b0000000000000000;
    rom[2894] = 16'b0001111111110000;
    rom[2895] = 16'b0001111111110000;
    rom[2896] = 16'b0000000001100000;
    rom[2897] = 16'b0000000011000000;
    rom[2898] = 16'b0000000011000000;
    rom[2899] = 16'b0000000110000000;
    rom[2900] = 16'b0000001100000000;
    rom[2901] = 16'b0000011000000000;
    rom[2902] = 16'b0000011000000000;
    rom[2903] = 16'b0000110000000000;
    rom[2904] = 16'b0001111111110000;
    rom[2905] = 16'b0001111111110000;
    rom[2906] = 16'b0000000000000000;
    rom[2907] = 16'b0000000000000000;
    rom[2908] = 16'b0000000000000000;
    rom[2909] = 16'b0000000000000000;
    rom[2910] = 16'b0000000000000000;
    rom[2911] = 16'b0000000000000000;

    // ASCII 123 (91): '{'
    rom[2912] = 16'b0000000000000000;
    rom[2913] = 16'b0000000000000000;
    rom[2914] = 16'b0000000000000000;
    rom[2915] = 16'b0000000000000000;
    rom[2916] = 16'b0000000011100000;
    rom[2917] = 16'b0000000111100000;
    rom[2918] = 16'b0000001110000000;
    rom[2919] = 16'b0000001100000000;
    rom[2920] = 16'b0000001100000000;
    rom[2921] = 16'b0000001100000000;
    rom[2922] = 16'b0000001100000000;
    rom[2923] = 16'b0000001100000000;
    rom[2924] = 16'b0000011100000000;
    rom[2925] = 16'b0001111000000000;
    rom[2926] = 16'b0001111000000000;
    rom[2927] = 16'b0000011100000000;
    rom[2928] = 16'b0000001100000000;
    rom[2929] = 16'b0000001100000000;
    rom[2930] = 16'b0000001100000000;
    rom[2931] = 16'b0000001100000000;
    rom[2932] = 16'b0000001100000000;
    rom[2933] = 16'b0000001100000000;
    rom[2934] = 16'b0000001100000000;
    rom[2935] = 16'b0000001110000000;
    rom[2936] = 16'b0000000111100000;
    rom[2937] = 16'b0000000011100000;
    rom[2938] = 16'b0000000000000000;
    rom[2939] = 16'b0000000000000000;
    rom[2940] = 16'b0000000000000000;
    rom[2941] = 16'b0000000000000000;
    rom[2942] = 16'b0000000000000000;
    rom[2943] = 16'b0000000000000000;

    // ASCII 124 (92): '|'
    rom[2944] = 16'b0000000000000000;
    rom[2945] = 16'b0000000110000000;
    rom[2946] = 16'b0000000110000000;
    rom[2947] = 16'b0000000110000000;
    rom[2948] = 16'b0000000110000000;
    rom[2949] = 16'b0000000110000000;
    rom[2950] = 16'b0000000110000000;
    rom[2951] = 16'b0000000110000000;
    rom[2952] = 16'b0000000110000000;
    rom[2953] = 16'b0000000110000000;
    rom[2954] = 16'b0000000110000000;
    rom[2955] = 16'b0000000110000000;
    rom[2956] = 16'b0000000110000000;
    rom[2957] = 16'b0000000110000000;
    rom[2958] = 16'b0000000110000000;
    rom[2959] = 16'b0000000110000000;
    rom[2960] = 16'b0000000110000000;
    rom[2961] = 16'b0000000110000000;
    rom[2962] = 16'b0000000110000000;
    rom[2963] = 16'b0000000110000000;
    rom[2964] = 16'b0000000110000000;
    rom[2965] = 16'b0000000110000000;
    rom[2966] = 16'b0000000110000000;
    rom[2967] = 16'b0000000110000000;
    rom[2968] = 16'b0000000110000000;
    rom[2969] = 16'b0000000000000000;
    rom[2970] = 16'b0000000000000000;
    rom[2971] = 16'b0000000000000000;
    rom[2972] = 16'b0000000000000000;
    rom[2973] = 16'b0000000000000000;
    rom[2974] = 16'b0000000000000000;
    rom[2975] = 16'b0000000000000000;

    // ASCII 125 (93): '}'
    rom[2976] = 16'b0000000000000000;
    rom[2977] = 16'b0000000000000000;
    rom[2978] = 16'b0000000000000000;
    rom[2979] = 16'b0000000000000000;
    rom[2980] = 16'b0000111000000000;
    rom[2981] = 16'b0000111100000000;
    rom[2982] = 16'b0000001110000000;
    rom[2983] = 16'b0000000110000000;
    rom[2984] = 16'b0000000110000000;
    rom[2985] = 16'b0000000110000000;
    rom[2986] = 16'b0000000110000000;
    rom[2987] = 16'b0000000110000000;
    rom[2988] = 16'b0000000111000000;
    rom[2989] = 16'b0000000011110000;
    rom[2990] = 16'b0000000011110000;
    rom[2991] = 16'b0000000111000000;
    rom[2992] = 16'b0000000110000000;
    rom[2993] = 16'b0000000110000000;
    rom[2994] = 16'b0000000110000000;
    rom[2995] = 16'b0000000110000000;
    rom[2996] = 16'b0000000110000000;
    rom[2997] = 16'b0000000110000000;
    rom[2998] = 16'b0000000110000000;
    rom[2999] = 16'b0000001110000000;
    rom[3000] = 16'b0000111100000000;
    rom[3001] = 16'b0000111000000000;
    rom[3002] = 16'b0000000000000000;
    rom[3003] = 16'b0000000000000000;
    rom[3004] = 16'b0000000000000000;
    rom[3005] = 16'b0000000000000000;
    rom[3006] = 16'b0000000000000000;
    rom[3007] = 16'b0000000000000000;

    // ASCII 126 (94): '~'
    rom[3008] = 16'b0000000000000000;
    rom[3009] = 16'b0000000000000000;
    rom[3010] = 16'b0000000000000000;
    rom[3011] = 16'b0000000000000000;
    rom[3012] = 16'b0000000000000000;
    rom[3013] = 16'b0000000000000000;
    rom[3014] = 16'b0000000000000000;
    rom[3015] = 16'b0000000000000000;
    rom[3016] = 16'b0000000000000000;
    rom[3017] = 16'b0000000000000000;
    rom[3018] = 16'b0000000000000000;
    rom[3019] = 16'b0000000000000000;
    rom[3020] = 16'b0000000000000000;
    rom[3021] = 16'b0000000000000000;
    rom[3022] = 16'b0000000000000000;
    rom[3023] = 16'b0000000000000000;
    rom[3024] = 16'b0000000000000000;
    rom[3025] = 16'b0000000000000000;
    rom[3026] = 16'b0000111000000000;
    rom[3027] = 16'b0001111100001100;
    rom[3028] = 16'b0011000110001100;
    rom[3029] = 16'b0011000011111000;
    rom[3030] = 16'b0000000001110000;
    rom[3031] = 16'b0000000000000000;
    rom[3032] = 16'b0000000000000000;
    rom[3033] = 16'b0000000000000000;
    rom[3034] = 16'b0000000000000000;
    rom[3035] = 16'b0000000000000000;
    rom[3036] = 16'b0000000000000000;
    rom[3037] = 16'b0000000000000000;
    rom[3038] = 16'b0000000000000000;
    rom[3039] = 16'b0000000000000000;

end

//=============================================================================
// ROM读取逻辑 (带流水线)
//=============================================================================
reg [15:0] char_data_reg;
reg [11:0] rom_addr;

always @(posedge clk) begin
    // 计算地址: (char_code - 32) * 32 + char_row
    if (char_code >= 32 && char_code <= 126) begin
        rom_addr <= (char_code - 32) * 32 + {7'd0, char_row};
        char_data_reg <= rom[rom_addr];
    end else begin
        char_data_reg <= 16'h0000;  // 非法字符显示空白
    end
end

assign char_data = char_data_reg;

endmodule
