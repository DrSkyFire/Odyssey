//=============================================================================
// 文件名: key_debounce.v
// 描述: 按键消抖模块
// 功能: 消除按键抖动，输出单脉冲信号
//=============================================================================

module key_debounce (
    input  wire clk,
    input  wire rst_n,
    input  wire key_in,             // 按键输入（低有效）
    output reg  key_pulse           // 按键脉冲输出（高有效，单周期）
);

//=============================================================================
// 参数定义
//=============================================================================
localparam DEBOUNCE_TIME = 20'd1_000_000;   // 消抖时间 10ms @ 100MHz

//=============================================================================
// 信号定义
//=============================================================================
reg [19:0] cnt;
reg        key_sync_0, key_sync_1;
reg        key_state;

//=============================================================================
// 按键同步（两级寄存器）
//=============================================================================
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        key_sync_0 <= 1'b1;
        key_sync_1 <= 1'b1;
    end else begin
        key_sync_0 <= key_in;
        key_sync_1 <= key_sync_0;
    end
end

//=============================================================================
// 消抖计数器
//=============================================================================
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        cnt <= 20'd0;
    end else begin
        if (key_sync_1 != key_state)
            cnt <= cnt + 1'b1;
        else
            cnt <= 20'd0;
    end
end

//=============================================================================
// 按键状态更新
//=============================================================================
always @(posedge clk or negedge rst_n) begin
    if (!rst_n)
        key_state <= 1'b1;
    else if (cnt == DEBOUNCE_TIME)
        key_state <= key_sync_1;
end

//=============================================================================
// 边沿检测 - 生成单脉冲
//=============================================================================
reg key_state_d1;

always @(posedge clk or negedge rst_n) begin
    if (!rst_n)
        key_state_d1 <= 1'b1;
    else
        key_state_d1 <= key_state;
end

always @(posedge clk or negedge rst_n) begin
    if (!rst_n)
        key_pulse <= 1'b0;
    else
        key_pulse <= key_state_d1 & ~key_state;  // 下降沿检测
end

endmodule