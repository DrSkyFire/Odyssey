//=============================================================================
// 文件名: char_rom_16x32.v
// 描述: 16x32点阵字符ROM - 支持0-9数字及常用字符
// 美观的大字体设计，适合HDMI显示
//
// 字符编码映射表:
// 数字: 0-9 → 编码 0-9
// 符号: '.'(10), ':'(11), '%'(12)
// 大写字母: 'C'(12), 'F'(16), 'H'(18), 'N'(23), 'S'(29), 'T'(30), 'U'(32)
// 小写字母: 'a'(17), 'e'(15), 'i'(19), 'k'(21), 'n'(24), 'o'(25), 'q'(27), 'r'(28), 'u'(31), 'w'(33), 'z'(14)
// 特殊符号: ':'(44), '%'(37)
//
// AI波形类型名称映射:
// - "Sine" = S(29) + i(19) + n(24) + e(15)
// - "Squr" = S(29) + q(27) + u(31) + r(28)
// - "Tria" = T(30) + r(28) + i(19) + a(17)
// - "Saw"  = S(29) + a(17) + w(33)
// - "Nois" = N(23) + o(25) + i(19) + s(29) [使用小写s]
// - "Unkn" = U(32) + n(24) + k(21) + n(24)
//=============================================================================

module char_rom_16x32 (
    input  wire [5:0]   char_code,      // 字符编码
    input  wire [4:0]   row,            // 行号 (0-31)
    output reg  [15:0]  pixel_row       // 16位像素行数据
);

always @(*) begin
    case (char_code)
        //=====================================================
        // '0' - ASCII 48
        //=====================================================
        6'd0: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0001111111111000;
                5'd2:  pixel_row = 16'b0011111111111100;
                5'd3:  pixel_row = 16'b0111110000111110;
                5'd4:  pixel_row = 16'b0111100000011110;
                5'd5:  pixel_row = 16'b1111000000001111;
                5'd6:  pixel_row = 16'b1111000000001111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1110000000000111;
                5'd9:  pixel_row = 16'b1110000000000111;
                5'd10: pixel_row = 16'b1110000000000111;
                5'd11: pixel_row = 16'b1110000000000111;
                5'd12: pixel_row = 16'b1110000000000111;
                5'd13: pixel_row = 16'b1110000000000111;
                5'd14: pixel_row = 16'b1110000000000111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                5'd17: pixel_row = 16'b1110000000000111;
                5'd18: pixel_row = 16'b1110000000000111;
                5'd19: pixel_row = 16'b1110000000000111;
                5'd20: pixel_row = 16'b1110000000000111;
                5'd21: pixel_row = 16'b1110000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1110000000000111;
                5'd24: pixel_row = 16'b1111000000001111;
                5'd25: pixel_row = 16'b1111000000001111;
                5'd26: pixel_row = 16'b0111100000011110;
                5'd27: pixel_row = 16'b0111110000111110;
                5'd28: pixel_row = 16'b0011111111111100;
                5'd29: pixel_row = 16'b0001111111111000;
                5'd30: pixel_row = 16'b0000111111110000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '1' - ASCII 49
        //=====================================================
        6'd1: begin
            case (row)
                5'd0:  pixel_row = 16'b0000001110000000;
                5'd1:  pixel_row = 16'b0000011110000000;
                5'd2:  pixel_row = 16'b0000111110000000;
                5'd3:  pixel_row = 16'b0001111110000000;
                5'd4:  pixel_row = 16'b0011111110000000;
                5'd5:  pixel_row = 16'b0011100110000000;
                5'd6:  pixel_row = 16'b0000000110000000;
                5'd7:  pixel_row = 16'b0000000110000000;
                5'd8:  pixel_row = 16'b0000000110000000;
                5'd9:  pixel_row = 16'b0000000110000000;
                5'd10: pixel_row = 16'b0000000110000000;
                5'd11: pixel_row = 16'b0000000110000000;
                5'd12: pixel_row = 16'b0000000110000000;
                5'd13: pixel_row = 16'b0000000110000000;
                5'd14: pixel_row = 16'b0000000110000000;
                5'd15: pixel_row = 16'b0000000110000000;
                5'd16: pixel_row = 16'b0000000110000000;
                5'd17: pixel_row = 16'b0000000110000000;
                5'd18: pixel_row = 16'b0000000110000000;
                5'd19: pixel_row = 16'b0000000110000000;
                5'd20: pixel_row = 16'b0000000110000000;
                5'd21: pixel_row = 16'b0000000110000000;
                5'd22: pixel_row = 16'b0000000110000000;
                5'd23: pixel_row = 16'b0000000110000000;
                5'd24: pixel_row = 16'b0000000110000000;
                5'd25: pixel_row = 16'b0000000110000000;
                5'd26: pixel_row = 16'b0000000110000000;
                5'd27: pixel_row = 16'b0111111111111110;
                5'd28: pixel_row = 16'b0111111111111110;
                5'd29: pixel_row = 16'b0111111111111110;
                5'd30: pixel_row = 16'b0111111111111110;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '2' - ASCII 50
        //=====================================================
        6'd2: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0011111111111100;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111100000011110;
                5'd4:  pixel_row = 16'b1110000000001111;
                5'd5:  pixel_row = 16'b1110000000000111;
                5'd6:  pixel_row = 16'b0000000000000111;
                5'd7:  pixel_row = 16'b0000000000000111;
                5'd8:  pixel_row = 16'b0000000000001111;
                5'd9:  pixel_row = 16'b0000000000011110;
                5'd10: pixel_row = 16'b0000000000111100;
                5'd11: pixel_row = 16'b0000000001111000;
                5'd12: pixel_row = 16'b0000000011110000;
                5'd13: pixel_row = 16'b0000000111100000;
                5'd14: pixel_row = 16'b0000001111000000;
                5'd15: pixel_row = 16'b0000011110000000;
                5'd16: pixel_row = 16'b0000111100000000;
                5'd17: pixel_row = 16'b0001111000000000;
                5'd18: pixel_row = 16'b0011110000000000;
                5'd19: pixel_row = 16'b0111100000000000;
                5'd20: pixel_row = 16'b0111000000000000;
                5'd21: pixel_row = 16'b1110000000000000;
                5'd22: pixel_row = 16'b1110000000000000;
                5'd23: pixel_row = 16'b1110000000000000;
                5'd24: pixel_row = 16'b1110000000000000;
                5'd25: pixel_row = 16'b1111000000000000;
                5'd26: pixel_row = 16'b1111111111111111;
                5'd27: pixel_row = 16'b1111111111111111;
                5'd28: pixel_row = 16'b1111111111111111;
                5'd29: pixel_row = 16'b1111111111111111;
                5'd30: pixel_row = 16'b1111111111111111;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '3' - ASCII 51
        //=====================================================
        6'd3: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0011111111111100;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111000000011110;
                5'd4:  pixel_row = 16'b1110000000001111;
                5'd5:  pixel_row = 16'b0000000000000111;
                5'd6:  pixel_row = 16'b0000000000000111;
                5'd7:  pixel_row = 16'b0000000000001110;
                5'd8:  pixel_row = 16'b0000000000111100;
                5'd9:  pixel_row = 16'b0000000111111000;
                5'd10: pixel_row = 16'b0000000111111000;
                5'd11: pixel_row = 16'b0000000111111000;
                5'd12: pixel_row = 16'b0000000111111000;
                5'd13: pixel_row = 16'b0000000111111000;
                5'd14: pixel_row = 16'b0000000000111100;
                5'd15: pixel_row = 16'b0000000000001110;
                5'd16: pixel_row = 16'b0000000000000111;
                5'd17: pixel_row = 16'b0000000000000111;
                5'd18: pixel_row = 16'b0000000000000111;
                5'd19: pixel_row = 16'b0000000000000111;
                5'd20: pixel_row = 16'b0000000000000111;
                5'd21: pixel_row = 16'b0000000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1110000000001111;
                5'd24: pixel_row = 16'b1111000000001111;
                5'd25: pixel_row = 16'b0111100000011110;
                5'd26: pixel_row = 16'b0111110000111110;
                5'd27: pixel_row = 16'b0011111111111100;
                5'd28: pixel_row = 16'b0001111111111000;
                5'd29: pixel_row = 16'b0000111111110000;
                5'd30: pixel_row = 16'b0000011111100000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '4' - ASCII 52
        //=====================================================
        6'd4: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000001111000;
                5'd1:  pixel_row = 16'b0000000011111000;
                5'd2:  pixel_row = 16'b0000000111111000;
                5'd3:  pixel_row = 16'b0000000111011000;
                5'd4:  pixel_row = 16'b0000001110011000;
                5'd5:  pixel_row = 16'b0000011100011000;
                5'd6:  pixel_row = 16'b0000011100011000;
                5'd7:  pixel_row = 16'b0000111000011000;
                5'd8:  pixel_row = 16'b0001110000011000;
                5'd9:  pixel_row = 16'b0011100000011000;
                5'd10: pixel_row = 16'b0011100000011000;
                5'd11: pixel_row = 16'b0111000000011000;
                5'd12: pixel_row = 16'b1110000000011000;
                5'd13: pixel_row = 16'b1110000000011000;
                5'd14: pixel_row = 16'b1100000000011000;
                5'd15: pixel_row = 16'b1111111111111111;
                5'd16: pixel_row = 16'b1111111111111111;
                5'd17: pixel_row = 16'b1111111111111111;
                5'd18: pixel_row = 16'b0000000000011000;
                5'd19: pixel_row = 16'b0000000000011000;
                5'd20: pixel_row = 16'b0000000000011000;
                5'd21: pixel_row = 16'b0000000000011000;
                5'd22: pixel_row = 16'b0000000000011000;
                5'd23: pixel_row = 16'b0000000000011000;
                5'd24: pixel_row = 16'b0000000000011000;
                5'd25: pixel_row = 16'b0000000000011000;
                5'd26: pixel_row = 16'b0000000000011000;
                5'd27: pixel_row = 16'b0000000000011000;
                5'd28: pixel_row = 16'b0000000000011000;
                5'd29: pixel_row = 16'b0000000000011000;
                5'd30: pixel_row = 16'b0000000000011000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '5' - ASCII 53
        //=====================================================
        6'd5: begin
            case (row)
                5'd0:  pixel_row = 16'b0111111111111110;
                5'd1:  pixel_row = 16'b0111111111111110;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111000000000000;
                5'd4:  pixel_row = 16'b0111000000000000;
                5'd5:  pixel_row = 16'b1110000000000000;
                5'd6:  pixel_row = 16'b1110000000000000;
                5'd7:  pixel_row = 16'b1110000000000000;
                5'd8:  pixel_row = 16'b1110111111100000;
                5'd9:  pixel_row = 16'b1111111111111000;
                5'd10: pixel_row = 16'b1111111111111100;
                5'd11: pixel_row = 16'b1111100000111110;
                5'd12: pixel_row = 16'b1110000000011110;
                5'd13: pixel_row = 16'b0000000000001111;
                5'd14: pixel_row = 16'b0000000000000111;
                5'd15: pixel_row = 16'b0000000000000111;
                5'd16: pixel_row = 16'b0000000000000111;
                5'd17: pixel_row = 16'b0000000000000111;
                5'd18: pixel_row = 16'b0000000000000111;
                5'd19: pixel_row = 16'b0000000000000111;
                5'd20: pixel_row = 16'b0000000000000111;
                5'd21: pixel_row = 16'b0000000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1110000000001111;
                5'd24: pixel_row = 16'b1111000000001111;
                5'd25: pixel_row = 16'b0111100000011110;
                5'd26: pixel_row = 16'b0111110000111110;
                5'd27: pixel_row = 16'b0011111111111100;
                5'd28: pixel_row = 16'b0001111111111000;
                5'd29: pixel_row = 16'b0000111111110000;
                5'd30: pixel_row = 16'b0000011111100000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '6' - ASCII 54
        //=====================================================
        6'd6: begin
            case (row)
                5'd0:  pixel_row = 16'b0000011111110000;
                5'd1:  pixel_row = 16'b0001111111111000;
                5'd2:  pixel_row = 16'b0011111111111100;
                5'd3:  pixel_row = 16'b0111110000000000;
                5'd4:  pixel_row = 16'b0111100000000000;
                5'd5:  pixel_row = 16'b1111000000000000;
                5'd6:  pixel_row = 16'b1110000000000000;
                5'd7:  pixel_row = 16'b1110000000000000;
                5'd8:  pixel_row = 16'b1110011111100000;
                5'd9:  pixel_row = 16'b1110111111111000;
                5'd10: pixel_row = 16'b1111111111111100;
                5'd11: pixel_row = 16'b1111110000111110;
                5'd12: pixel_row = 16'b1111100000011110;
                5'd13: pixel_row = 16'b1111000000001111;
                5'd14: pixel_row = 16'b1110000000000111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                5'd17: pixel_row = 16'b1110000000000111;
                5'd18: pixel_row = 16'b1110000000000111;
                5'd19: pixel_row = 16'b1110000000000111;
                5'd20: pixel_row = 16'b1110000000000111;
                5'd21: pixel_row = 16'b1110000000000111;
                5'd22: pixel_row = 16'b1110000000001111;
                5'd23: pixel_row = 16'b1111000000001111;
                5'd24: pixel_row = 16'b0111100000011110;
                5'd25: pixel_row = 16'b0111110000111110;
                5'd26: pixel_row = 16'b0011111111111100;
                5'd27: pixel_row = 16'b0001111111111000;
                5'd28: pixel_row = 16'b0000111111110000;
                5'd29: pixel_row = 16'b0000011111100000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '7' - ASCII 55
        //=====================================================
        6'd7: begin
            case (row)
                5'd0:  pixel_row = 16'b1111111111111111;
                5'd1:  pixel_row = 16'b1111111111111111;
                5'd2:  pixel_row = 16'b1111111111111111;
                5'd3:  pixel_row = 16'b1111111111111111;
                5'd4:  pixel_row = 16'b0000000000000111;
                5'd5:  pixel_row = 16'b0000000000001110;
                5'd6:  pixel_row = 16'b0000000000011100;
                5'd7:  pixel_row = 16'b0000000000111000;
                5'd8:  pixel_row = 16'b0000000000111000;
                5'd9:  pixel_row = 16'b0000000001110000;
                5'd10: pixel_row = 16'b0000000011100000;
                5'd11: pixel_row = 16'b0000000011100000;
                5'd12: pixel_row = 16'b0000000111000000;
                5'd13: pixel_row = 16'b0000000111000000;
                5'd14: pixel_row = 16'b0000001110000000;
                5'd15: pixel_row = 16'b0000001110000000;
                5'd16: pixel_row = 16'b0000011100000000;
                5'd17: pixel_row = 16'b0000011100000000;
                5'd18: pixel_row = 16'b0000111000000000;
                5'd19: pixel_row = 16'b0000111000000000;
                5'd20: pixel_row = 16'b0001110000000000;
                5'd21: pixel_row = 16'b0001110000000000;
                5'd22: pixel_row = 16'b0011100000000000;
                5'd23: pixel_row = 16'b0011100000000000;
                5'd24: pixel_row = 16'b0111000000000000;
                5'd25: pixel_row = 16'b0111000000000000;
                5'd26: pixel_row = 16'b1110000000000000;
                5'd27: pixel_row = 16'b1110000000000000;
                5'd28: pixel_row = 16'b1110000000000000;
                5'd29: pixel_row = 16'b1100000000000000;
                5'd30: pixel_row = 16'b1100000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '8' - ASCII 56
        //=====================================================
        6'd8: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0011111111111100;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111100000011110;
                5'd4:  pixel_row = 16'b1111000000001111;
                5'd5:  pixel_row = 16'b1110000000000111;
                5'd6:  pixel_row = 16'b1110000000000111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1111000000001111;
                5'd9:  pixel_row = 16'b0111100000011110;
                5'd10: pixel_row = 16'b0011111111111100;
                5'd11: pixel_row = 16'b0001111111111000;
                5'd12: pixel_row = 16'b0011111111111100;
                5'd13: pixel_row = 16'b0111100000011110;
                5'd14: pixel_row = 16'b1111000000001111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                5'd17: pixel_row = 16'b1110000000000111;
                5'd18: pixel_row = 16'b1110000000000111;
                5'd19: pixel_row = 16'b1110000000000111;
                5'd20: pixel_row = 16'b1110000000000111;
                5'd21: pixel_row = 16'b1110000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1111000000001111;
                5'd24: pixel_row = 16'b0111100000011110;
                5'd25: pixel_row = 16'b0111110000111110;
                5'd26: pixel_row = 16'b0011111111111100;
                5'd27: pixel_row = 16'b0001111111111000;
                5'd28: pixel_row = 16'b0000111111110000;
                5'd29: pixel_row = 16'b0000011111100000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '9' - ASCII 57
        //=====================================================
        6'd9: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0011111111111100;
                5'd2:  pixel_row = 16'b0111111111111110;
                5'd3:  pixel_row = 16'b0111110000111110;
                5'd4:  pixel_row = 16'b1111100000011111;
                5'd5:  pixel_row = 16'b1111000000001111;
                5'd6:  pixel_row = 16'b1110000000000111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1110000000000111;
                5'd9:  pixel_row = 16'b1110000000000111;
                5'd10: pixel_row = 16'b1110000000000111;
                5'd11: pixel_row = 16'b1110000000000111;
                5'd12: pixel_row = 16'b1110000000000111;
                5'd13: pixel_row = 16'b1111000000000111;
                5'd14: pixel_row = 16'b1111100000001111;
                5'd15: pixel_row = 16'b0111110000011111;
                5'd16: pixel_row = 16'b0111111111111111;
                5'd17: pixel_row = 16'b0011111111110111;
                5'd18: pixel_row = 16'b0001111110000111;
                5'd19: pixel_row = 16'b0000000000000111;
                5'd20: pixel_row = 16'b0000000000000111;
                5'd21: pixel_row = 16'b0000000000001111;
                5'd22: pixel_row = 16'b0000000000001110;
                5'd23: pixel_row = 16'b0000000000011110;
                5'd24: pixel_row = 16'b0000000000111100;
                5'd25: pixel_row = 16'b0000000001111000;
                5'd26: pixel_row = 16'b0111110011110000;
                5'd27: pixel_row = 16'b0111111111100000;
                5'd28: pixel_row = 16'b0011111111000000;
                5'd29: pixel_row = 16'b0001111110000000;
                5'd30: pixel_row = 16'b0000111100000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '.' - 点号 (ASCII 46)
        //=====================================================
        6'd10: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000000000000000;
                5'd5:  pixel_row = 16'b0000000000000000;
                5'd6:  pixel_row = 16'b0000000000000000;
                5'd7:  pixel_row = 16'b0000000000000000;
                5'd8:  pixel_row = 16'b0000000000000000;
                5'd9:  pixel_row = 16'b0000000000000000;
                5'd10: pixel_row = 16'b0000000000000000;
                5'd11: pixel_row = 16'b0000000000000000;
                5'd12: pixel_row = 16'b0000000000000000;
                5'd13: pixel_row = 16'b0000000000000000;
                5'd14: pixel_row = 16'b0000000000000000;
                5'd15: pixel_row = 16'b0000000000000000;
                5'd16: pixel_row = 16'b0000000000000000;
                5'd17: pixel_row = 16'b0000000000000000;
                5'd18: pixel_row = 16'b0000000000000000;
                5'd19: pixel_row = 16'b0000000000000000;
                5'd20: pixel_row = 16'b0000000000000000;
                5'd21: pixel_row = 16'b0000000000000000;
                5'd22: pixel_row = 16'b0000000000000000;
                5'd23: pixel_row = 16'b0000000000000000;
                5'd24: pixel_row = 16'b0000011111000000;
                5'd25: pixel_row = 16'b0000011111000000;
                5'd26: pixel_row = 16'b0000011111000000;
                5'd27: pixel_row = 16'b0000011111000000;
                5'd28: pixel_row = 16'b0000011111000000;
                5'd29: pixel_row = 16'b0000011111000000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // ':' - 冒号 (ASCII 58)
        //=====================================================
        6'd11: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000000000000000;
                5'd5:  pixel_row = 16'b0000000000000000;
                5'd6:  pixel_row = 16'b0000000000000000;
                5'd7:  pixel_row = 16'b0000011111000000;
                5'd8:  pixel_row = 16'b0000011111000000;
                5'd9:  pixel_row = 16'b0000011111000000;
                5'd10: pixel_row = 16'b0000011111000000;
                5'd11: pixel_row = 16'b0000011111000000;
                5'd12: pixel_row = 16'b0000011111000000;
                5'd13: pixel_row = 16'b0000000000000000;
                5'd14: pixel_row = 16'b0000000000000000;
                5'd15: pixel_row = 16'b0000000000000000;
                5'd16: pixel_row = 16'b0000000000000000;
                5'd17: pixel_row = 16'b0000000000000000;
                5'd18: pixel_row = 16'b0000000000000000;
                5'd19: pixel_row = 16'b0000011111000000;
                5'd20: pixel_row = 16'b0000011111000000;
                5'd21: pixel_row = 16'b0000011111000000;
                5'd22: pixel_row = 16'b0000011111000000;
                5'd23: pixel_row = 16'b0000011111000000;
                5'd24: pixel_row = 16'b0000011111000000;
                5'd25: pixel_row = 16'b0000000000000000;
                5'd26: pixel_row = 16'b0000000000000000;
                5'd27: pixel_row = 16'b0000000000000000;
                5'd28: pixel_row = 16'b0000000000000000;
                5'd29: pixel_row = 16'b0000000000000000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '%' - 百分号 (ASCII 37)
        //=====================================================
        6'd12: begin
            case (row)
                5'd0:  pixel_row = 16'b0111000000000110;
                5'd1:  pixel_row = 16'b1101100000001110;
                5'd2:  pixel_row = 16'b1101100000011100;
                5'd3:  pixel_row = 16'b1101100000111000;
                5'd4:  pixel_row = 16'b1101100000110000;
                5'd5:  pixel_row = 16'b0111000001110000;
                5'd6:  pixel_row = 16'b0000000011100000;
                5'd7:  pixel_row = 16'b0000000111000000;
                5'd8:  pixel_row = 16'b0000000110000000;
                5'd9:  pixel_row = 16'b0000001110000000;
                5'd10: pixel_row = 16'b0000011100000000;
                5'd11: pixel_row = 16'b0000011000000000;
                5'd12: pixel_row = 16'b0000111000000000;
                5'd13: pixel_row = 16'b0000110000000000;
                5'd14: pixel_row = 16'b0001110000000000;
                5'd15: pixel_row = 16'b0011100000000000;
                5'd16: pixel_row = 16'b0011000000000000;
                5'd17: pixel_row = 16'b0111000000000000;
                5'd18: pixel_row = 16'b0110000000111000;
                5'd19: pixel_row = 16'b1110000001101100;
                5'd20: pixel_row = 16'b1100000001101100;
                5'd21: pixel_row = 16'b1100000001101100;
                5'd22: pixel_row = 16'b0000000001101100;
                5'd23: pixel_row = 16'b0000000000111000;
                5'd24: pixel_row = 16'b0000000000000000;
                5'd25: pixel_row = 16'b0000000000000000;
                5'd26: pixel_row = 16'b0000000000000000;
                5'd27: pixel_row = 16'b0000000000000000;
                5'd28: pixel_row = 16'b0000000000000000;
                5'd29: pixel_row = 16'b0000000000000000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'H' - 字母H (ASCII 72)
        //=====================================================
        6'd13: begin
            case (row)
                5'd0:  pixel_row = 16'b1110000000000111;
                5'd1:  pixel_row = 16'b1110000000000111;
                5'd2:  pixel_row = 16'b1110000000000111;
                5'd3:  pixel_row = 16'b1110000000000111;
                5'd4:  pixel_row = 16'b1110000000000111;
                5'd5:  pixel_row = 16'b1110000000000111;
                5'd6:  pixel_row = 16'b1110000000000111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1110000000000111;
                5'd9:  pixel_row = 16'b1110000000000111;
                5'd10: pixel_row = 16'b1110000000000111;
                5'd11: pixel_row = 16'b1111111111111111;
                5'd12: pixel_row = 16'b1111111111111111;
                5'd13: pixel_row = 16'b1111111111111111;
                5'd14: pixel_row = 16'b1111111111111111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                5'd17: pixel_row = 16'b1110000000000111;
                5'd18: pixel_row = 16'b1110000000000111;
                5'd19: pixel_row = 16'b1110000000000111;
                5'd20: pixel_row = 16'b1110000000000111;
                5'd21: pixel_row = 16'b1110000000000111;
                5'd22: pixel_row = 16'b1110000000000111;
                5'd23: pixel_row = 16'b1110000000000111;
                5'd24: pixel_row = 16'b1110000000000111;
                5'd25: pixel_row = 16'b1110000000000111;
                5'd26: pixel_row = 16'b1110000000000111;
                5'd27: pixel_row = 16'b1110000000000111;
                5'd28: pixel_row = 16'b1110000000000111;
                5'd29: pixel_row = 16'b1110000000000111;
                5'd30: pixel_row = 16'b1110000000000111;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'z' - 字母z (ASCII 122)
        //=====================================================
        6'd14: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000000000000000;
                5'd5:  pixel_row = 16'b0111111111111110;
                5'd6:  pixel_row = 16'b0111111111111110;
                5'd7:  pixel_row = 16'b0111111111111110;
                5'd8:  pixel_row = 16'b0000000000111110;
                5'd9:  pixel_row = 16'b0000000001111100;
                5'd10: pixel_row = 16'b0000000011111000;
                5'd11: pixel_row = 16'b0000000111110000;
                5'd12: pixel_row = 16'b0000001111100000;
                5'd13: pixel_row = 16'b0000011111000000;
                5'd14: pixel_row = 16'b0000111110000000;
                5'd15: pixel_row = 16'b0001111100000000;
                5'd16: pixel_row = 16'b0011111000000000;
                5'd17: pixel_row = 16'b0111110000000000;
                5'd18: pixel_row = 16'b0111100000000000;
                5'd19: pixel_row = 16'b1111000000000000;
                5'd20: pixel_row = 16'b1110000000000000;
                5'd21: pixel_row = 16'b1111111111111110;
                5'd22: pixel_row = 16'b1111111111111110;
                5'd23: pixel_row = 16'b1111111111111110;
                5'd24: pixel_row = 16'b0000000000000000;
                5'd25: pixel_row = 16'b0000000000000000;
                5'd26: pixel_row = 16'b0000000000000000;
                5'd27: pixel_row = 16'b0000000000000000;
                5'd28: pixel_row = 16'b0000000000000000;
                5'd29: pixel_row = 16'b0000000000000000;
                5'd30: pixel_row = 16'b0000000000000000;
                5'd31: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'e' - 字母e (编码15)
        //=====================================================
        6'd15: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000111111100000;
                5'd5:  pixel_row = 16'b0011111111110000;
                5'd6:  pixel_row = 16'b0111100001111000;
                5'd7:  pixel_row = 16'b1110000000111100;
                5'd8:  pixel_row = 16'b1110000000111100;
                5'd9:  pixel_row = 16'b1111111111111100;
                5'd10: pixel_row = 16'b1111111111111100;
                5'd11: pixel_row = 16'b1111111111111100;
                5'd12: pixel_row = 16'b1110000000000000;
                5'd13: pixel_row = 16'b1110000000000000;
                5'd14: pixel_row = 16'b1110000000111100;
                5'd15: pixel_row = 16'b0111100001111000;
                5'd16: pixel_row = 16'b0011111111110000;
                5'd17: pixel_row = 16'b0000111111100000;
                5'd18: pixel_row = 16'b0000000000000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'a' - 字母a (编码17)
        //=====================================================
        6'd17: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000111111100000;
                5'd5:  pixel_row = 16'b0011111111110000;
                5'd6:  pixel_row = 16'b0111100001111000;
                5'd7:  pixel_row = 16'b0000000000111100;
                5'd8:  pixel_row = 16'b0000111111111100;
                5'd9:  pixel_row = 16'b0111111111111100;
                5'd10: pixel_row = 16'b1111000000111100;
                5'd11: pixel_row = 16'b1110000000111100;
                5'd12: pixel_row = 16'b1110000000111100;
                5'd13: pixel_row = 16'b1111000001111100;
                5'd14: pixel_row = 16'b0111111111111100;
                5'd15: pixel_row = 16'b0011111110111100;
                5'd16: pixel_row = 16'b0000000000000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'i' - 字母i (编码19)
        //=====================================================
        6'd19: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000011100000000;
                5'd2:  pixel_row = 16'b0000011100000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0001111100000000;
                5'd5:  pixel_row = 16'b0001111100000000;
                5'd6:  pixel_row = 16'b0000011100000000;
                5'd7:  pixel_row = 16'b0000011100000000;
                5'd8:  pixel_row = 16'b0000011100000000;
                5'd9:  pixel_row = 16'b0000011100000000;
                5'd10: pixel_row = 16'b0000011100000000;
                5'd11: pixel_row = 16'b0000011100000000;
                5'd12: pixel_row = 16'b0000011100000000;
                5'd13: pixel_row = 16'b0000011100000000;
                5'd14: pixel_row = 16'b0000011100000000;
                5'd15: pixel_row = 16'b0001111111000000;
                5'd16: pixel_row = 16'b0001111111000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'n' - 字母n (编码24)
        //=====================================================
        6'd24: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b1110111110000000;
                5'd5:  pixel_row = 16'b1111111111000000;
                5'd6:  pixel_row = 16'b1111000111100000;
                5'd7:  pixel_row = 16'b1110000011100000;
                5'd8:  pixel_row = 16'b1110000011100000;
                5'd9:  pixel_row = 16'b1110000011100000;
                5'd10: pixel_row = 16'b1110000011100000;
                5'd11: pixel_row = 16'b1110000011100000;
                5'd12: pixel_row = 16'b1110000011100000;
                5'd13: pixel_row = 16'b1110000011100000;
                5'd14: pixel_row = 16'b1110000011100000;
                5'd15: pixel_row = 16'b1110000011100000;
                5'd16: pixel_row = 16'b1110000011100000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'o' - 字母o (编码25)
        //=====================================================
        6'd25: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000111111000000;
                5'd5:  pixel_row = 16'b0011111111110000;
                5'd6:  pixel_row = 16'b0111000001111000;
                5'd7:  pixel_row = 16'b1110000000111000;
                5'd8:  pixel_row = 16'b1110000000111000;
                5'd9:  pixel_row = 16'b1110000000111000;
                5'd10: pixel_row = 16'b1110000000111000;
                5'd11: pixel_row = 16'b1110000000111000;
                5'd12: pixel_row = 16'b0111000001111000;
                5'd13: pixel_row = 16'b0011111111110000;
                5'd14: pixel_row = 16'b0000111111000000;
                5'd15: pixel_row = 16'b0000000000000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'S' - 字母S (编码29)
        //=====================================================
        6'd29: begin
            case (row)
                5'd0:  pixel_row = 16'b0000111111110000;
                5'd1:  pixel_row = 16'b0011111111111100;
                5'd2:  pixel_row = 16'b0111100000111110;
                5'd3:  pixel_row = 16'b1110000000011110;
                5'd4:  pixel_row = 16'b1110000000000000;
                5'd5:  pixel_row = 16'b1111000000000000;
                5'd6:  pixel_row = 16'b0111100000000000;
                5'd7:  pixel_row = 16'b0011111110000000;
                5'd8:  pixel_row = 16'b0001111111110000;
                5'd9:  pixel_row = 16'b0000011111111000;
                5'd10: pixel_row = 16'b0000000111111100;
                5'd11: pixel_row = 16'b0000000001111100;
                5'd12: pixel_row = 16'b0000000000111100;
                5'd13: pixel_row = 16'b0000000000111100;
                5'd14: pixel_row = 16'b1110000000111100;
                5'd15: pixel_row = 16'b1111000001111000;
                5'd16: pixel_row = 16'b0111111111110000;
                5'd17: pixel_row = 16'b0001111111100000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'C' - 字母C (编码12) - 修正已存在的，改为字母C而非数字
        //=====================================================
        6'd12: begin
            case (row)
                5'd0:  pixel_row = 16'b0000011111110000;
                5'd1:  pixel_row = 16'b0001111111111000;
                5'd2:  pixel_row = 16'b0011111111111100;
                5'd3:  pixel_row = 16'b0111100000111110;
                5'd4:  pixel_row = 16'b1110000000011110;
                5'd5:  pixel_row = 16'b1110000000000000;
                5'd6:  pixel_row = 16'b1110000000000000;
                5'd7:  pixel_row = 16'b1110000000000000;
                5'd8:  pixel_row = 16'b1110000000000000;
                5'd9:  pixel_row = 16'b1110000000000000;
                5'd10: pixel_row = 16'b1110000000000000;
                5'd11: pixel_row = 16'b1110000000000000;
                5'd12: pixel_row = 16'b1110000000000000;
                5'd13: pixel_row = 16'b1110000000000000;
                5'd14: pixel_row = 16'b1110000000000000;
                5'd15: pixel_row = 16'b1110000000000000;
                5'd16: pixel_row = 16'b1110000000000000;
                5'd17: pixel_row = 16'b1110000000011110;
                5'd18: pixel_row = 16'b0111100000111110;
                5'd19: pixel_row = 16'b0011111111111100;
                5'd20: pixel_row = 16'b0001111111111000;
                5'd21: pixel_row = 16'b0000011111110000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'H' - 字母H (编码18) - 修正编码18为字母H
        //=====================================================
        6'd18: begin
            case (row)
                5'd0:  pixel_row = 16'b1110000000000111;
                5'd1:  pixel_row = 16'b1110000000000111;
                5'd2:  pixel_row = 16'b1110000000000111;
                5'd3:  pixel_row = 16'b1110000000000111;
                5'd4:  pixel_row = 16'b1110000000000111;
                5'd5:  pixel_row = 16'b1110000000000111;
                5'd6:  pixel_row = 16'b1110000000000111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1111111111111111;
                5'd9:  pixel_row = 16'b1111111111111111;
                5'd10: pixel_row = 16'b1111111111111111;
                5'd11: pixel_row = 16'b1110000000000111;
                5'd12: pixel_row = 16'b1110000000000111;
                5'd13: pixel_row = 16'b1110000000000111;
                5'd14: pixel_row = 16'b1110000000000111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                5'd17: pixel_row = 16'b1110000000000111;
                5'd18: pixel_row = 16'b1110000000000111;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'q' - 字母q (编码27)
        //=====================================================
        6'd27: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000111110111000;
                5'd4:  pixel_row = 16'b0011111111111100;
                5'd5:  pixel_row = 16'b0111000001111100;
                5'd6:  pixel_row = 16'b1110000000111100;
                5'd7:  pixel_row = 16'b1110000000111100;
                5'd8:  pixel_row = 16'b1110000000111100;
                5'd9:  pixel_row = 16'b0111000001111100;
                5'd10: pixel_row = 16'b0011111111111100;
                5'd11: pixel_row = 16'b0000111110111100;
                5'd12: pixel_row = 16'b0000000000111100;
                5'd13: pixel_row = 16'b0000000000111100;
                5'd14: pixel_row = 16'b0000000000111100;
                5'd15: pixel_row = 16'b0000000000111100;
                5'd16: pixel_row = 16'b0000000000111100;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'r' - 字母r (编码28)
        //=====================================================
        6'd28: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b1110011111000000;
                5'd5:  pixel_row = 16'b1110111111100000;
                5'd6:  pixel_row = 16'b1111110001110000;
                5'd7:  pixel_row = 16'b1111100000000000;
                5'd8:  pixel_row = 16'b1111000000000000;
                5'd9:  pixel_row = 16'b1110000000000000;
                5'd10: pixel_row = 16'b1110000000000000;
                5'd11: pixel_row = 16'b1110000000000000;
                5'd12: pixel_row = 16'b1110000000000000;
                5'd13: pixel_row = 16'b1110000000000000;
                5'd14: pixel_row = 16'b1110000000000000;
                5'd15: pixel_row = 16'b1110000000000000;
                5'd16: pixel_row = 16'b1110000000000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'T' - 字母T (编码30)
        //=====================================================
        6'd30: begin
            case (row)
                5'd0:  pixel_row = 16'b1111111111111111;
                5'd1:  pixel_row = 16'b1111111111111111;
                5'd2:  pixel_row = 16'b1111111111111111;
                5'd3:  pixel_row = 16'b0000001110000000;
                5'd4:  pixel_row = 16'b0000001110000000;
                5'd5:  pixel_row = 16'b0000001110000000;
                5'd6:  pixel_row = 16'b0000001110000000;
                5'd7:  pixel_row = 16'b0000001110000000;
                5'd8:  pixel_row = 16'b0000001110000000;
                5'd9:  pixel_row = 16'b0000001110000000;
                5'd10: pixel_row = 16'b0000001110000000;
                5'd11: pixel_row = 16'b0000001110000000;
                5'd12: pixel_row = 16'b0000001110000000;
                5'd13: pixel_row = 16'b0000001110000000;
                5'd14: pixel_row = 16'b0000001110000000;
                5'd15: pixel_row = 16'b0000001110000000;
                5'd16: pixel_row = 16'b0000001110000000;
                5'd17: pixel_row = 16'b0000001110000000;
                5'd18: pixel_row = 16'b0000001110000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'u' - 字母u (编码31)
        //=====================================================
        6'd31: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b1110000000111000;
                5'd5:  pixel_row = 16'b1110000000111000;
                5'd6:  pixel_row = 16'b1110000000111000;
                5'd7:  pixel_row = 16'b1110000000111000;
                5'd8:  pixel_row = 16'b1110000000111000;
                5'd9:  pixel_row = 16'b1110000000111000;
                5'd10: pixel_row = 16'b1110000000111000;
                5'd11: pixel_row = 16'b1110000000111000;
                5'd12: pixel_row = 16'b1110000000111000;
                5'd13: pixel_row = 16'b1111000001111000;
                5'd14: pixel_row = 16'b0111111111111000;
                5'd15: pixel_row = 16'b0011111110111000;
                5'd16: pixel_row = 16'b0000000000000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'w' - 字母w (编码33)
        //=====================================================
        6'd33: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b1110000000001110;
                5'd5:  pixel_row = 16'b1110000000001110;
                5'd6:  pixel_row = 16'b1110000000001110;
                5'd7:  pixel_row = 16'b1110000000001110;
                5'd8:  pixel_row = 16'b1110000111001110;
                5'd9:  pixel_row = 16'b1110001111101110;
                5'd10: pixel_row = 16'b1110011101111110;
                5'd11: pixel_row = 16'b1110111000011110;
                5'd12: pixel_row = 16'b1111110000111100;
                5'd13: pixel_row = 16'b0111100000111000;
                5'd14: pixel_row = 16'b0111000000110000;
                5'd15: pixel_row = 16'b0000000000000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'k' - 字母k (编码21)
        //=====================================================
        6'd21: begin
            case (row)
                5'd0:  pixel_row = 16'b1110000000000000;
                5'd1:  pixel_row = 16'b1110000000000000;
                5'd2:  pixel_row = 16'b1110000000000000;
                5'd3:  pixel_row = 16'b1110000000000000;
                5'd4:  pixel_row = 16'b1110000001111000;
                5'd5:  pixel_row = 16'b1110000011110000;
                5'd6:  pixel_row = 16'b1110000111100000;
                5'd7:  pixel_row = 16'b1110001111000000;
                5'd8:  pixel_row = 16'b1110011110000000;
                5'd9:  pixel_row = 16'b1110111100000000;
                5'd10: pixel_row = 16'b1111111000000000;
                5'd11: pixel_row = 16'b1111011100000000;
                5'd12: pixel_row = 16'b1110001111000000;
                5'd13: pixel_row = 16'b1110000111100000;
                5'd14: pixel_row = 16'b1110000011110000;
                5'd15: pixel_row = 16'b1110000001111000;
                5'd16: pixel_row = 16'b1110000000111100;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'U' - 字母U (编码32) - 大写U
        //=====================================================
        6'd32: begin
            case (row)
                5'd0:  pixel_row = 16'b1110000000000111;
                5'd1:  pixel_row = 16'b1110000000000111;
                5'd2:  pixel_row = 16'b1110000000000111;
                5'd3:  pixel_row = 16'b1110000000000111;
                5'd4:  pixel_row = 16'b1110000000000111;
                5'd5:  pixel_row = 16'b1110000000000111;
                5'd6:  pixel_row = 16'b1110000000000111;
                5'd7:  pixel_row = 16'b1110000000000111;
                5'd8:  pixel_row = 16'b1110000000000111;
                5'd9:  pixel_row = 16'b1110000000000111;
                5'd10: pixel_row = 16'b1110000000000111;
                5'd11: pixel_row = 16'b1110000000000111;
                5'd12: pixel_row = 16'b1110000000000111;
                5'd13: pixel_row = 16'b1111000000001111;
                5'd14: pixel_row = 16'b0111100000011110;
                5'd15: pixel_row = 16'b0011111111111100;
                5'd16: pixel_row = 16'b0001111111111000;
                5'd17: pixel_row = 16'b0000111111110000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'N' - 字母N (编码23) - 大写N
        //=====================================================
        6'd23: begin
            case (row)
                5'd0:  pixel_row = 16'b1110000000000111;
                5'd1:  pixel_row = 16'b1111000000000111;
                5'd2:  pixel_row = 16'b1111100000000111;
                5'd3:  pixel_row = 16'b1111110000000111;
                5'd4:  pixel_row = 16'b1111111000000111;
                5'd5:  pixel_row = 16'b1110111100000111;
                5'd6:  pixel_row = 16'b1110011110000111;
                5'd7:  pixel_row = 16'b1110001111000111;
                5'd8:  pixel_row = 16'b1110000111100111;
                5'd9:  pixel_row = 16'b1110000011110111;
                5'd10: pixel_row = 16'b1110000001111111;
                5'd11: pixel_row = 16'b1110000000111111;
                5'd12: pixel_row = 16'b1110000000011111;
                5'd13: pixel_row = 16'b1110000000001111;
                5'd14: pixel_row = 16'b1110000000000111;
                5'd15: pixel_row = 16'b1110000000000111;
                5'd16: pixel_row = 16'b1110000000000111;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // ':' - 冒号 (编码44)
        //=====================================================
        6'd44: begin
            case (row)
                5'd0:  pixel_row = 16'b0000000000000000;
                5'd1:  pixel_row = 16'b0000000000000000;
                5'd2:  pixel_row = 16'b0000000000000000;
                5'd3:  pixel_row = 16'b0000000000000000;
                5'd4:  pixel_row = 16'b0000011100000000;
                5'd5:  pixel_row = 16'b0000111110000000;
                5'd6:  pixel_row = 16'b0000111110000000;
                5'd7:  pixel_row = 16'b0000011100000000;
                5'd8:  pixel_row = 16'b0000000000000000;
                5'd9:  pixel_row = 16'b0000000000000000;
                5'd10: pixel_row = 16'b0000000000000000;
                5'd11: pixel_row = 16'b0000000000000000;
                5'd12: pixel_row = 16'b0000000000000000;
                5'd13: pixel_row = 16'b0000011100000000;
                5'd14: pixel_row = 16'b0000111110000000;
                5'd15: pixel_row = 16'b0000111110000000;
                5'd16: pixel_row = 16'b0000011100000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // '%' - 百分号 (编码37)
        //=====================================================
        6'd37: begin
            case (row)
                5'd0:  pixel_row = 16'b0111000000000110;
                5'd1:  pixel_row = 16'b1101100000001110;
                5'd2:  pixel_row = 16'b1101100000011100;
                5'd3:  pixel_row = 16'b1101100000111000;
                5'd4:  pixel_row = 16'b1101100000110000;
                5'd5:  pixel_row = 16'b0111000001110000;
                5'd6:  pixel_row = 16'b0000000011100000;
                5'd7:  pixel_row = 16'b0000000111000000;
                5'd8:  pixel_row = 16'b0000000110000000;
                5'd9:  pixel_row = 16'b0000001110000000;
                5'd10: pixel_row = 16'b0000011100000000;
                5'd11: pixel_row = 16'b0000011000000000;
                5'd12: pixel_row = 16'b0000111000000000;
                5'd13: pixel_row = 16'b0000110000000000;
                5'd14: pixel_row = 16'b0001110000000000;
                5'd15: pixel_row = 16'b0011100000111000;
                5'd16: pixel_row = 16'b0011000001101100;
                5'd17: pixel_row = 16'b0111000001101100;
                5'd18: pixel_row = 16'b0110000001101100;
                5'd19: pixel_row = 16'b1110000001101100;
                5'd20: pixel_row = 16'b1100000000111000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 'F' - 字母F (编码16) - 用于"Freq"
        //=====================================================
        6'd16: begin
            case (row)
                5'd0:  pixel_row = 16'b1111111111111110;
                5'd1:  pixel_row = 16'b1111111111111110;
                5'd2:  pixel_row = 16'b1111111111111110;
                5'd3:  pixel_row = 16'b1110000000000000;
                5'd4:  pixel_row = 16'b1110000000000000;
                5'd5:  pixel_row = 16'b1110000000000000;
                5'd6:  pixel_row = 16'b1110000000000000;
                5'd7:  pixel_row = 16'b1111111111110000;
                5'd8:  pixel_row = 16'b1111111111110000;
                5'd9:  pixel_row = 16'b1111111111110000;
                5'd10: pixel_row = 16'b1110000000000000;
                5'd11: pixel_row = 16'b1110000000000000;
                5'd12: pixel_row = 16'b1110000000000000;
                5'd13: pixel_row = 16'b1110000000000000;
                5'd14: pixel_row = 16'b1110000000000000;
                5'd15: pixel_row = 16'b1110000000000000;
                5'd16: pixel_row = 16'b1110000000000000;
                5'd17: pixel_row = 16'b1110000000000000;
                default: pixel_row = 16'b0000000000000000;
            endcase
        end
        
        //=====================================================
        // 空格 (ASCII 32) 和其他未定义字符
        //=====================================================
        default: pixel_row = 16'b0000000000000000;
    endcase
end

endmodule
