//=============================================================================
// 文件名称: ascii_rom_16x32.v
// 模块名称: ascii_rom_16x32
// 功能描述: 16×32像素ASCII字符ROM (支持ASCII码32-126)
//          包含: 数字0-9, 大小写字母A-Z/a-z, 常用符号
// 设计者  : AI Assistant
// 创建日期: 2025-10-26
//=============================================================================

module ascii_rom_16x32 (
    input        clk,
    input  [7:0] char_code,   // ASCII码 (32-126有效)
    input  [4:0] char_row,    // 字符行号 (0-31)
    output [15:0] char_data   // 16位字符行数据
);

//=============================================================================
// 字符ROM存储器
//=============================================================================
// ASCII 32-126 共95个字符, 每个字符32行×16位 = 512字节
// 总ROM大小: 95 × 512 = 47.5KB

reg [15:0] char_rom [0:3039];  // 95个字符 × 32行 = 3040行

//=============================================================================
// ROM初始化 (可选使用 $readmemh 从文件读取)
//=============================================================================
initial begin
    // 这里我们手动初始化常用字符
    // 您也可以使用: $readmemh("ascii_font_16x32.hex", char_rom);
    
    // 初始化所有字符为空白
    integer i;
    for (i = 0; i < 3040; i = i + 1) begin
        char_rom[i] = 16'h0000;
    end
    
    // ========== 空格 (ASCII 32 = 0) ==========
    // 保持全0
    
    // ========== ! (ASCII 33 = 1) ==========
    char_rom[1*32 + 8]  = 16'b0000001100000000;
    char_rom[1*32 + 9]  = 16'b0000001100000000;
    char_rom[1*32 + 10] = 16'b0000001100000000;
    char_rom[1*32 + 11] = 16'b0000001100000000;
    char_rom[1*32 + 12] = 16'b0000001100000000;
    char_rom[1*32 + 13] = 16'b0000001100000000;
    char_rom[1*32 + 14] = 16'b0000001100000000;
    char_rom[1*32 + 15] = 16'b0000001100000000;
    char_rom[1*32 + 16] = 16'b0000001100000000;
    char_rom[1*32 + 17] = 16'b0000001100000000;
    char_rom[1*32 + 18] = 16'b0000000000000000;
    char_rom[1*32 + 19] = 16'b0000000000000000;
    char_rom[1*32 + 20] = 16'b0000001100000000;
    char_rom[1*32 + 21] = 16'b0000001100000000;
    
    // ========== % (ASCII 37 = 5) ==========
    char_rom[5*32 + 8]  = 16'b0001100000011000;
    char_rom[5*32 + 9]  = 16'b0011110000110000;
    char_rom[5*32 + 10] = 16'b0011110000110000;
    char_rom[5*32 + 11] = 16'b0001100001100000;
    char_rom[5*32 + 12] = 16'b0000000001100000;
    char_rom[5*32 + 13] = 16'b0000000011000000;
    char_rom[5*32 + 14] = 16'b0000000011000000;
    char_rom[5*32 + 15] = 16'b0000000110000000;
    char_rom[5*32 + 16] = 16'b0000001100000000;
    char_rom[5*32 + 17] = 16'b0000001100000000;
    char_rom[5*32 + 18] = 16'b0000011000000000;
    char_rom[5*32 + 19] = 16'b0000110001100000;
    char_rom[5*32 + 20] = 16'b0000110011110000;
    char_rom[5*32 + 21] = 16'b0001100011110000;
    char_rom[5*32 + 22] = 16'b0001100001100000;
    
    // ========== . (ASCII 46 = 14) ==========
    char_rom[14*32 + 20] = 16'b0000011000000000;
    char_rom[14*32 + 21] = 16'b0000011000000000;
    
    // ========== : (ASCII 58 = 26) ==========
    char_rom[26*32 + 12] = 16'b0000011000000000;
    char_rom[26*32 + 13] = 16'b0000011000000000;
    char_rom[26*32 + 14] = 16'b0000000000000000;
    char_rom[26*32 + 15] = 16'b0000000000000000;
    char_rom[26*32 + 16] = 16'b0000000000000000;
    char_rom[26*32 + 17] = 16'b0000000000000000;
    char_rom[26*32 + 18] = 16'b0000011000000000;
    char_rom[26*32 + 19] = 16'b0000011000000000;
    
    // ========== 数字 0-9 (ASCII 48-57 = index 16-25) ==========
    
    // 0 (ASCII 48 = 16)
    char_rom[16*32 + 8]  = 16'b0000111111000000;
    char_rom[16*32 + 9]  = 16'b0011111111110000;
    char_rom[16*32 + 10] = 16'b0011000000110000;
    char_rom[16*32 + 11] = 16'b0011000000110000;
    char_rom[16*32 + 12] = 16'b0011000000110000;
    char_rom[16*32 + 13] = 16'b0011000000110000;
    char_rom[16*32 + 14] = 16'b0011000000110000;
    char_rom[16*32 + 15] = 16'b0011000000110000;
    char_rom[16*32 + 16] = 16'b0011000000110000;
    char_rom[16*32 + 17] = 16'b0011000000110000;
    char_rom[16*32 + 18] = 16'b0011000000110000;
    char_rom[16*32 + 19] = 16'b0011000000110000;
    char_rom[16*32 + 20] = 16'b0011111111110000;
    char_rom[16*32 + 21] = 16'b0000111111000000;
    
    // 1 (ASCII 49 = 17)
    char_rom[17*32 + 8]  = 16'b0000001100000000;
    char_rom[17*32 + 9]  = 16'b0000111100000000;
    char_rom[17*32 + 10] = 16'b0000001100000000;
    char_rom[17*32 + 11] = 16'b0000001100000000;
    char_rom[17*32 + 12] = 16'b0000001100000000;
    char_rom[17*32 + 13] = 16'b0000001100000000;
    char_rom[17*32 + 14] = 16'b0000001100000000;
    char_rom[17*32 + 15] = 16'b0000001100000000;
    char_rom[17*32 + 16] = 16'b0000001100000000;
    char_rom[17*32 + 17] = 16'b0000001100000000;
    char_rom[17*32 + 18] = 16'b0000001100000000;
    char_rom[17*32 + 19] = 16'b0000001100000000;
    char_rom[17*32 + 20] = 16'b0011111111110000;
    char_rom[17*32 + 21] = 16'b0011111111110000;
    
    // 2 (ASCII 50 = 18)
    char_rom[18*32 + 8]  = 16'b0000111111000000;
    char_rom[18*32 + 9]  = 16'b0011111111110000;
    char_rom[18*32 + 10] = 16'b0011000000110000;
    char_rom[18*32 + 11] = 16'b0000000000110000;
    char_rom[18*32 + 12] = 16'b0000000000110000;
    char_rom[18*32 + 13] = 16'b0000000001100000;
    char_rom[18*32 + 14] = 16'b0000000011000000;
    char_rom[18*32 + 15] = 16'b0000000110000000;
    char_rom[18*32 + 16] = 16'b0000001100000000;
    char_rom[18*32 + 17] = 16'b0000011000000000;
    char_rom[18*32 + 18] = 16'b0000110000000000;
    char_rom[18*32 + 19] = 16'b0011000000000000;
    char_rom[18*32 + 20] = 16'b0011111111110000;
    char_rom[18*32 + 21] = 16'b0011111111110000;
    
    // 3 (ASCII 51 = 19)
    char_rom[19*32 + 8]  = 16'b0000111111000000;
    char_rom[19*32 + 9]  = 16'b0011111111110000;
    char_rom[19*32 + 10] = 16'b0011000000110000;
    char_rom[19*32 + 11] = 16'b0000000000110000;
    char_rom[19*32 + 12] = 16'b0000000000110000;
    char_rom[19*32 + 13] = 16'b0000001111110000;
    char_rom[19*32 + 14] = 16'b0000001111110000;
    char_rom[19*32 + 15] = 16'b0000000000110000;
    char_rom[19*32 + 16] = 16'b0000000000110000;
    char_rom[19*32 + 17] = 16'b0000000000110000;
    char_rom[19*32 + 18] = 16'b0000000000110000;
    char_rom[19*32 + 19] = 16'b0011000000110000;
    char_rom[19*32 + 20] = 16'b0011111111110000;
    char_rom[19*32 + 21] = 16'b0000111111000000;
    
    // 4 (ASCII 52 = 20)
    char_rom[20*32 + 8]  = 16'b0000000011000000;
    char_rom[20*32 + 9]  = 16'b0000000111000000;
    char_rom[20*32 + 10] = 16'b0000001111000000;
    char_rom[20*32 + 11] = 16'b0000011011000000;
    char_rom[20*32 + 12] = 16'b0000110011000000;
    char_rom[20*32 + 13] = 16'b0001100011000000;
    char_rom[20*32 + 14] = 16'b0011000011000000;
    char_rom[20*32 + 15] = 16'b0011111111111000;
    char_rom[20*32 + 16] = 16'b0011111111111000;
    char_rom[20*32 + 17] = 16'b0000000011000000;
    char_rom[20*32 + 18] = 16'b0000000011000000;
    char_rom[20*32 + 19] = 16'b0000000011000000;
    char_rom[20*32 + 20] = 16'b0000000011000000;
    char_rom[20*32 + 21] = 16'b0000000011000000;
    
    // 5 (ASCII 53 = 21)
    char_rom[21*32 + 8]  = 16'b0011111111110000;
    char_rom[21*32 + 9]  = 16'b0011111111110000;
    char_rom[21*32 + 10] = 16'b0011000000000000;
    char_rom[21*32 + 11] = 16'b0011000000000000;
    char_rom[21*32 + 12] = 16'b0011000000000000;
    char_rom[21*32 + 13] = 16'b0011111111000000;
    char_rom[21*32 + 14] = 16'b0011111111110000;
    char_rom[21*32 + 15] = 16'b0000000000110000;
    char_rom[21*32 + 16] = 16'b0000000000110000;
    char_rom[21*32 + 17] = 16'b0000000000110000;
    char_rom[21*32 + 18] = 16'b0000000000110000;
    char_rom[21*32 + 19] = 16'b0011000000110000;
    char_rom[21*32 + 20] = 16'b0011111111110000;
    char_rom[21*32 + 21] = 16'b0000111111000000;
    
    // 6 (ASCII 54 = 22)
    char_rom[22*32 + 8]  = 16'b0000111111000000;
    char_rom[22*32 + 9]  = 16'b0011111111110000;
    char_rom[22*32 + 10] = 16'b0011000000110000;
    char_rom[22*32 + 11] = 16'b0011000000000000;
    char_rom[22*32 + 12] = 16'b0011000000000000;
    char_rom[22*32 + 13] = 16'b0011111111000000;
    char_rom[22*32 + 14] = 16'b0011111111110000;
    char_rom[22*32 + 15] = 16'b0011000000110000;
    char_rom[22*32 + 16] = 16'b0011000000110000;
    char_rom[22*32 + 17] = 16'b0011000000110000;
    char_rom[22*32 + 18] = 16'b0011000000110000;
    char_rom[22*32 + 19] = 16'b0011000000110000;
    char_rom[22*32 + 20] = 16'b0011111111110000;
    char_rom[22*32 + 21] = 16'b0000111111000000;
    
    // 7 (ASCII 55 = 23)
    char_rom[23*32 + 8]  = 16'b0011111111110000;
    char_rom[23*32 + 9]  = 16'b0011111111110000;
    char_rom[23*32 + 10] = 16'b0000000000110000;
    char_rom[23*32 + 11] = 16'b0000000000110000;
    char_rom[23*32 + 12] = 16'b0000000001100000;
    char_rom[23*32 + 13] = 16'b0000000011000000;
    char_rom[23*32 + 14] = 16'b0000000110000000;
    char_rom[23*32 + 15] = 16'b0000001100000000;
    char_rom[23*32 + 16] = 16'b0000011000000000;
    char_rom[23*32 + 17] = 16'b0000110000000000;
    char_rom[23*32 + 18] = 16'b0001100000000000;
    char_rom[23*32 + 19] = 16'b0001100000000000;
    char_rom[23*32 + 20] = 16'b0001100000000000;
    char_rom[23*32 + 21] = 16'b0001100000000000;
    
    // 8 (ASCII 56 = 24)
    char_rom[24*32 + 8]  = 16'b0000111111000000;
    char_rom[24*32 + 9]  = 16'b0011111111110000;
    char_rom[24*32 + 10] = 16'b0011000000110000;
    char_rom[24*32 + 11] = 16'b0011000000110000;
    char_rom[24*32 + 12] = 16'b0011000000110000;
    char_rom[24*32 + 13] = 16'b0000111111000000;
    char_rom[24*32 + 14] = 16'b0000111111000000;
    char_rom[24*32 + 15] = 16'b0011000000110000;
    char_rom[24*32 + 16] = 16'b0011000000110000;
    char_rom[24*32 + 17] = 16'b0011000000110000;
    char_rom[24*32 + 18] = 16'b0011000000110000;
    char_rom[24*32 + 19] = 16'b0011000000110000;
    char_rom[24*32 + 20] = 16'b0011111111110000;
    char_rom[24*32 + 21] = 16'b0000111111000000;
    
    // 9 (ASCII 57 = 25)
    char_rom[25*32 + 8]  = 16'b0000111111000000;
    char_rom[25*32 + 9]  = 16'b0011111111110000;
    char_rom[25*32 + 10] = 16'b0011000000110000;
    char_rom[25*32 + 11] = 16'b0011000000110000;
    char_rom[25*32 + 12] = 16'b0011000000110000;
    char_rom[25*32 + 13] = 16'b0011111111110000;
    char_rom[25*32 + 14] = 16'b0000111111110000;
    char_rom[25*32 + 15] = 16'b0000000000110000;
    char_rom[25*32 + 16] = 16'b0000000000110000;
    char_rom[25*32 + 17] = 16'b0000000000110000;
    char_rom[25*32 + 18] = 16'b0000000000110000;
    char_rom[25*32 + 19] = 16'b0011000000110000;
    char_rom[25*32 + 20] = 16'b0011111111110000;
    char_rom[25*32 + 21] = 16'b0000111111000000;
    
    // ========== 大写字母 A-Z (ASCII 65-90 = index 33-58) ==========
    
    // A (ASCII 65 = 33)
    char_rom[33*32 + 8]  = 16'b0000011110000000;
    char_rom[33*32 + 9]  = 16'b0000111111000000;
    char_rom[33*32 + 10] = 16'b0001100001100000;
    char_rom[33*32 + 11] = 16'b0011000000110000;
    char_rom[33*32 + 12] = 16'b0011000000110000;
    char_rom[33*32 + 13] = 16'b0011000000110000;
    char_rom[33*32 + 14] = 16'b0011111111110000;
    char_rom[33*32 + 15] = 16'b0011111111110000;
    char_rom[33*32 + 16] = 16'b0011000000110000;
    char_rom[33*32 + 17] = 16'b0011000000110000;
    char_rom[33*32 + 18] = 16'b0011000000110000;
    char_rom[33*32 + 19] = 16'b0011000000110000;
    char_rom[33*32 + 20] = 16'b0011000000110000;
    char_rom[33*32 + 21] = 16'b0011000000110000;
    
    // C (ASCII 67 = 35)
    char_rom[35*32 + 8]  = 16'b0000111111000000;
    char_rom[35*32 + 9]  = 16'b0011111111110000;
    char_rom[35*32 + 10] = 16'b0011000000110000;
    char_rom[35*32 + 11] = 16'b0011000000000000;
    char_rom[35*32 + 12] = 16'b0011000000000000;
    char_rom[35*32 + 13] = 16'b0011000000000000;
    char_rom[35*32 + 14] = 16'b0011000000000000;
    char_rom[35*32 + 15] = 16'b0011000000000000;
    char_rom[35*32 + 16] = 16'b0011000000000000;
    char_rom[35*32 + 17] = 16'b0011000000000000;
    char_rom[35*32 + 18] = 16'b0011000000000000;
    char_rom[35*32 + 19] = 16'b0011000000110000;
    char_rom[35*32 + 20] = 16'b0011111111110000;
    char_rom[35*32 + 21] = 16'b0000111111000000;
    
    // D (ASCII 68 = 36)
    char_rom[36*32 + 8]  = 16'b0011111110000000;
    char_rom[36*32 + 9]  = 16'b0011111111100000;
    char_rom[36*32 + 10] = 16'b0011000001110000;
    char_rom[36*32 + 11] = 16'b0011000000110000;
    char_rom[36*32 + 12] = 16'b0011000000110000;
    char_rom[36*32 + 13] = 16'b0011000000110000;
    char_rom[36*32 + 14] = 16'b0011000000110000;
    char_rom[36*32 + 15] = 16'b0011000000110000;
    char_rom[36*32 + 16] = 16'b0011000000110000;
    char_rom[36*32 + 17] = 16'b0011000000110000;
    char_rom[36*32 + 18] = 16'b0011000001110000;
    char_rom[36*32 + 19] = 16'b0011111111100000;
    char_rom[36*32 + 20] = 16'b0011111110000000;
    
    // F (ASCII 70 = 38)
    char_rom[38*32 + 8]  = 16'b0011111111110000;
    char_rom[38*32 + 9]  = 16'b0011111111110000;
    char_rom[38*32 + 10] = 16'b0011000000000000;
    char_rom[38*32 + 11] = 16'b0011000000000000;
    char_rom[38*32 + 12] = 16'b0011000000000000;
    char_rom[38*32 + 13] = 16'b0011111111000000;
    char_rom[38*32 + 14] = 16'b0011111111000000;
    char_rom[38*32 + 15] = 16'b0011000000000000;
    char_rom[38*32 + 16] = 16'b0011000000000000;
    char_rom[38*32 + 17] = 16'b0011000000000000;
    char_rom[38*32 + 18] = 16'b0011000000000000;
    char_rom[38*32 + 19] = 16'b0011000000000000;
    char_rom[38*32 + 20] = 16'b0011000000000000;
    char_rom[38*32 + 21] = 16'b0011000000000000;
    
    // H (ASCII 72 = 40)
    char_rom[40*32 + 8]  = 16'b0011000000110000;
    char_rom[40*32 + 9]  = 16'b0011000000110000;
    char_rom[40*32 + 10] = 16'b0011000000110000;
    char_rom[40*32 + 11] = 16'b0011000000110000;
    char_rom[40*32 + 12] = 16'b0011000000110000;
    char_rom[40*32 + 13] = 16'b0011111111110000;
    char_rom[40*32 + 14] = 16'b0011111111110000;
    char_rom[40*32 + 15] = 16'b0011000000110000;
    char_rom[40*32 + 16] = 16'b0011000000110000;
    char_rom[40*32 + 17] = 16'b0011000000110000;
    char_rom[40*32 + 18] = 16'b0011000000110000;
    char_rom[40*32 + 19] = 16'b0011000000110000;
    char_rom[40*32 + 20] = 16'b0011000000110000;
    char_rom[40*32 + 21] = 16'b0011000000110000;
    
    // P (ASCII 80 = 48)
    char_rom[48*32 + 8]  = 16'b0011111111000000;
    char_rom[48*32 + 9]  = 16'b0011111111110000;
    char_rom[48*32 + 10] = 16'b0011000000110000;
    char_rom[48*32 + 11] = 16'b0011000000110000;
    char_rom[48*32 + 12] = 16'b0011000000110000;
    char_rom[48*32 + 13] = 16'b0011111111110000;
    char_rom[48*32 + 14] = 16'b0011111111000000;
    char_rom[48*32 + 15] = 16'b0011000000000000;
    char_rom[48*32 + 16] = 16'b0011000000000000;
    char_rom[48*32 + 17] = 16'b0011000000000000;
    char_rom[48*32 + 18] = 16'b0011000000000000;
    char_rom[48*32 + 19] = 16'b0011000000000000;
    char_rom[48*32 + 20] = 16'b0011000000000000;
    
    // S (ASCII 83 = 51)
    char_rom[51*32 + 8]  = 16'b0000111111000000;
    char_rom[51*32 + 9]  = 16'b0011111111110000;
    char_rom[51*32 + 10] = 16'b0011000000110000;
    char_rom[51*32 + 11] = 16'b0011000000000000;
    char_rom[51*32 + 12] = 16'b0011000000000000;
    char_rom[51*32 + 13] = 16'b0001111111000000;
    char_rom[51*32 + 14] = 16'b0000111111110000;
    char_rom[51*32 + 15] = 16'b0000000000110000;
    char_rom[51*32 + 16] = 16'b0000000000110000;
    char_rom[51*32 + 17] = 16'b0000000000110000;
    char_rom[51*32 + 18] = 16'b0000000000110000;
    char_rom[51*32 + 19] = 16'b0011000000110000;
    char_rom[51*32 + 20] = 16'b0011111111110000;
    char_rom[51*32 + 21] = 16'b0000111111000000;
    
    // T (ASCII 84 = 52)
    char_rom[52*32 + 8]  = 16'b0011111111110000;
    char_rom[52*32 + 9]  = 16'b0011111111110000;
    char_rom[52*32 + 10] = 16'b0000001100000000;
    char_rom[52*32 + 11] = 16'b0000001100000000;
    char_rom[52*32 + 12] = 16'b0000001100000000;
    char_rom[52*32 + 13] = 16'b0000001100000000;
    char_rom[52*32 + 14] = 16'b0000001100000000;
    char_rom[52*32 + 15] = 16'b0000001100000000;
    char_rom[52*32 + 16] = 16'b0000001100000000;
    char_rom[52*32 + 17] = 16'b0000001100000000;
    char_rom[52*32 + 18] = 16'b0000001100000000;
    char_rom[52*32 + 19] = 16'b0000001100000000;
    char_rom[52*32 + 20] = 16'b0000001100000000;
    char_rom[52*32 + 21] = 16'b0000001100000000;
    
    // 更多字母可以继续添加...
    // 为了简化,您可以使用字体生成工具创建完整字库
end

//=============================================================================
// 字符数据输出 (带流水线)
//=============================================================================
reg [15:0] char_data_reg;
reg [10:0] rom_addr;

always @(posedge clk) begin
    // 计算ROM地址: (char_code - 32) * 32 + char_row
    // ASCII 32-126 映射到 index 0-94
    if (char_code >= 32 && char_code <= 126) begin
        rom_addr <= (char_code - 32) * 32 + char_row;
    end else begin
        rom_addr <= 0;  // 非法字符显示为空格
    end
    
    // 读取字符数据
    char_data_reg <= char_rom[rom_addr];
end

assign char_data = char_data_reg;

endmodule
